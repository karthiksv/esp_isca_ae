`timescale 1ps / 1ps
module fft2_Mul_32Ux32U_32U_4(
          in2,
          in1,
          out1,
          clk,
          clr
);
   input [31:0] in2;
   input [31:0] in1;
   output [31:0] out1;
   input clk;
   input clr;
wire mul_22_8_n_0, mul_22_8_n_1, mul_22_8_n_2, mul_22_8_n_4, mul_22_8_n_5,
     mul_22_8_n_6, mul_22_8_n_8, mul_22_8_n_9, mul_22_8_n_10, mul_22_8_n_11,
     mul_22_8_n_12, mul_22_8_n_13, mul_22_8_n_14, mul_22_8_n_15, mul_22_8_n_16,
     mul_22_8_n_17, mul_22_8_n_18, mul_22_8_n_19, mul_22_8_n_20, mul_22_8_n_21,
     mul_22_8_n_22, mul_22_8_n_23, mul_22_8_n_24, mul_22_8_n_25, mul_22_8_n_26,
     mul_22_8_n_27, mul_22_8_n_29, mul_22_8_n_30, mul_22_8_n_31, mul_22_8_n_32,
     mul_22_8_n_33, mul_22_8_n_34, mul_22_8_n_35, mul_22_8_n_36, mul_22_8_n_37,
     mul_22_8_n_38, mul_22_8_n_39, mul_22_8_n_40, mul_22_8_n_41, mul_22_8_n_42,
     mul_22_8_n_43, mul_22_8_n_44, mul_22_8_n_45, mul_22_8_n_46, mul_22_8_n_48,
     mul_22_8_n_49, mul_22_8_n_50, mul_22_8_n_51, mul_22_8_n_52, mul_22_8_n_53,
     mul_22_8_n_54, mul_22_8_n_55, mul_22_8_n_56, mul_22_8_n_57, mul_22_8_n_58,
     mul_22_8_n_59, mul_22_8_n_60, mul_22_8_n_61, mul_22_8_n_62, mul_22_8_n_63,
     mul_22_8_n_64, mul_22_8_n_66, mul_22_8_n_67, mul_22_8_n_68, mul_22_8_n_69,
     mul_22_8_n_70, mul_22_8_n_71, mul_22_8_n_72, mul_22_8_n_73, mul_22_8_n_74,
     mul_22_8_n_75, mul_22_8_n_76, mul_22_8_n_77, mul_22_8_n_78, mul_22_8_n_79,
     mul_22_8_n_80, mul_22_8_n_81, mul_22_8_n_82, mul_22_8_n_83, mul_22_8_n_84,
     mul_22_8_n_85, mul_22_8_n_86, mul_22_8_n_87, mul_22_8_n_88, mul_22_8_n_89,
     mul_22_8_n_90, mul_22_8_n_91, mul_22_8_n_92, mul_22_8_n_93, mul_22_8_n_94,
     mul_22_8_n_95, mul_22_8_n_96, mul_22_8_n_97, mul_22_8_n_98, mul_22_8_n_99,
     mul_22_8_n_100, mul_22_8_n_101, mul_22_8_n_102, mul_22_8_n_103,
     mul_22_8_n_104, mul_22_8_n_105, mul_22_8_n_106, mul_22_8_n_107,
     mul_22_8_n_108, mul_22_8_n_109, mul_22_8_n_110, mul_22_8_n_111,
     mul_22_8_n_112, mul_22_8_n_113, mul_22_8_n_114, mul_22_8_n_115,
     mul_22_8_n_116, mul_22_8_n_117, mul_22_8_n_118, mul_22_8_n_119,
     mul_22_8_n_120, mul_22_8_n_121, mul_22_8_n_122, mul_22_8_n_123,
     mul_22_8_n_124, mul_22_8_n_125, mul_22_8_n_126, mul_22_8_n_127,
     mul_22_8_n_128, mul_22_8_n_129, mul_22_8_n_130, mul_22_8_n_131,
     mul_22_8_n_132, mul_22_8_n_133, mul_22_8_n_134, mul_22_8_n_135,
     mul_22_8_n_136, mul_22_8_n_137, mul_22_8_n_138, mul_22_8_n_139,
     mul_22_8_n_140, mul_22_8_n_141, mul_22_8_n_142, mul_22_8_n_143,
     mul_22_8_n_144, mul_22_8_n_145, mul_22_8_n_146, mul_22_8_n_147,
     mul_22_8_n_148, mul_22_8_n_149, mul_22_8_n_150, mul_22_8_n_151,
     mul_22_8_n_152, mul_22_8_n_153, mul_22_8_n_154, mul_22_8_n_155,
     mul_22_8_n_156, mul_22_8_n_157, mul_22_8_n_158, mul_22_8_n_159,
     mul_22_8_n_160, mul_22_8_n_161, mul_22_8_n_162, mul_22_8_n_163,
     mul_22_8_n_164, mul_22_8_n_165, mul_22_8_n_166, mul_22_8_n_167,
     mul_22_8_n_168, mul_22_8_n_169, mul_22_8_n_170, mul_22_8_n_171,
     mul_22_8_n_172, mul_22_8_n_173, mul_22_8_n_174, mul_22_8_n_175,
     mul_22_8_n_176, mul_22_8_n_177, mul_22_8_n_178, mul_22_8_n_179,
     mul_22_8_n_180, mul_22_8_n_181, mul_22_8_n_182, mul_22_8_n_183,
     mul_22_8_n_184, mul_22_8_n_185, mul_22_8_n_186, mul_22_8_n_187,
     mul_22_8_n_188, mul_22_8_n_189, mul_22_8_n_190, mul_22_8_n_191,
     mul_22_8_n_192, mul_22_8_n_193, mul_22_8_n_194, mul_22_8_n_195,
     mul_22_8_n_196, mul_22_8_n_197, mul_22_8_n_198, mul_22_8_n_199,
     mul_22_8_n_200, mul_22_8_n_201, mul_22_8_n_202, mul_22_8_n_203,
     mul_22_8_n_204, mul_22_8_n_205, mul_22_8_n_206, mul_22_8_n_207,
     mul_22_8_n_208, mul_22_8_n_209, mul_22_8_n_210, mul_22_8_n_211,
     mul_22_8_n_212, mul_22_8_n_213, mul_22_8_n_214, mul_22_8_n_215,
     mul_22_8_n_216, mul_22_8_n_217, mul_22_8_n_218, mul_22_8_n_219,
     mul_22_8_n_220, mul_22_8_n_221, mul_22_8_n_222, mul_22_8_n_223,
     mul_22_8_n_224, mul_22_8_n_225, mul_22_8_n_226, mul_22_8_n_227,
     mul_22_8_n_228, mul_22_8_n_229, mul_22_8_n_230, mul_22_8_n_231,
     mul_22_8_n_232, mul_22_8_n_233, mul_22_8_n_234, mul_22_8_n_235,
     mul_22_8_n_236, mul_22_8_n_237, mul_22_8_n_238, mul_22_8_n_239,
     mul_22_8_n_240, mul_22_8_n_241, mul_22_8_n_242, mul_22_8_n_244,
     mul_22_8_n_245, mul_22_8_n_246, mul_22_8_n_247, mul_22_8_n_248,
     mul_22_8_n_249, mul_22_8_n_250, mul_22_8_n_251, mul_22_8_n_252,
     mul_22_8_n_253, mul_22_8_n_254, mul_22_8_n_255, mul_22_8_n_256,
     mul_22_8_n_257, mul_22_8_n_258, mul_22_8_n_259, mul_22_8_n_260,
     mul_22_8_n_261, mul_22_8_n_262, mul_22_8_n_263, mul_22_8_n_264,
     mul_22_8_n_265, mul_22_8_n_266, mul_22_8_n_267, mul_22_8_n_268,
     mul_22_8_n_269, mul_22_8_n_270, mul_22_8_n_271, mul_22_8_n_272,
     mul_22_8_n_273, mul_22_8_n_274, mul_22_8_n_275, mul_22_8_n_276,
     mul_22_8_n_277, mul_22_8_n_278, mul_22_8_n_279, mul_22_8_n_280,
     mul_22_8_n_281, mul_22_8_n_282, mul_22_8_n_283, mul_22_8_n_284,
     mul_22_8_n_285, mul_22_8_n_286, mul_22_8_n_287, mul_22_8_n_288,
     mul_22_8_n_289, mul_22_8_n_290, mul_22_8_n_291, mul_22_8_n_292,
     mul_22_8_n_293, mul_22_8_n_294, mul_22_8_n_295, mul_22_8_n_296,
     mul_22_8_n_297, mul_22_8_n_298, mul_22_8_n_299, mul_22_8_n_300,
     mul_22_8_n_301, mul_22_8_n_302, mul_22_8_n_303, mul_22_8_n_304,
     mul_22_8_n_305, mul_22_8_n_306, mul_22_8_n_307, mul_22_8_n_308,
     mul_22_8_n_309, mul_22_8_n_310, mul_22_8_n_311, mul_22_8_n_312,
     mul_22_8_n_313, mul_22_8_n_314, mul_22_8_n_315, mul_22_8_n_316,
     mul_22_8_n_317, mul_22_8_n_318, mul_22_8_n_319, mul_22_8_n_320,
     mul_22_8_n_321, mul_22_8_n_322, mul_22_8_n_323, mul_22_8_n_324,
     mul_22_8_n_325, mul_22_8_n_326, mul_22_8_n_327, mul_22_8_n_328,
     mul_22_8_n_329, mul_22_8_n_330, mul_22_8_n_331, mul_22_8_n_332,
     mul_22_8_n_333, mul_22_8_n_334, mul_22_8_n_335, mul_22_8_n_336,
     mul_22_8_n_337, mul_22_8_n_338, mul_22_8_n_339, mul_22_8_n_340,
     mul_22_8_n_341, mul_22_8_n_342, mul_22_8_n_343, mul_22_8_n_344,
     mul_22_8_n_345, mul_22_8_n_346, mul_22_8_n_347, mul_22_8_n_348,
     mul_22_8_n_349, mul_22_8_n_350, mul_22_8_n_351, mul_22_8_n_352,
     mul_22_8_n_353, mul_22_8_n_354, mul_22_8_n_355, mul_22_8_n_356,
     mul_22_8_n_357, mul_22_8_n_358, mul_22_8_n_359, mul_22_8_n_360,
     mul_22_8_n_361, mul_22_8_n_362, mul_22_8_n_363, mul_22_8_n_364,
     mul_22_8_n_365, mul_22_8_n_366, mul_22_8_n_367, mul_22_8_n_368,
     mul_22_8_n_369, mul_22_8_n_370, mul_22_8_n_371, mul_22_8_n_372,
     mul_22_8_n_373, mul_22_8_n_374, mul_22_8_n_375, mul_22_8_n_376,
     mul_22_8_n_377, mul_22_8_n_378, mul_22_8_n_379, mul_22_8_n_380,
     mul_22_8_n_381, mul_22_8_n_382, mul_22_8_n_383, mul_22_8_n_384,
     mul_22_8_n_385, mul_22_8_n_386, mul_22_8_n_387, mul_22_8_n_388,
     mul_22_8_n_389, mul_22_8_n_390, mul_22_8_n_391, mul_22_8_n_392,
     mul_22_8_n_393, mul_22_8_n_394, mul_22_8_n_395, mul_22_8_n_396,
     mul_22_8_n_397, mul_22_8_n_398, mul_22_8_n_399, mul_22_8_n_400,
     mul_22_8_n_401, mul_22_8_n_402, mul_22_8_n_403, mul_22_8_n_404,
     mul_22_8_n_405, mul_22_8_n_406, mul_22_8_n_407, mul_22_8_n_408,
     mul_22_8_n_409, mul_22_8_n_410, mul_22_8_n_411, mul_22_8_n_412,
     mul_22_8_n_413, mul_22_8_n_414, mul_22_8_n_415, mul_22_8_n_416,
     mul_22_8_n_417, mul_22_8_n_418, mul_22_8_n_419, mul_22_8_n_420,
     mul_22_8_n_421, mul_22_8_n_422, mul_22_8_n_423, mul_22_8_n_424,
     mul_22_8_n_425, mul_22_8_n_426, mul_22_8_n_427, mul_22_8_n_428,
     mul_22_8_n_429, mul_22_8_n_430, mul_22_8_n_431, mul_22_8_n_432,
     mul_22_8_n_433, mul_22_8_n_434, mul_22_8_n_435, mul_22_8_n_436,
     mul_22_8_n_437, mul_22_8_n_438, mul_22_8_n_439, mul_22_8_n_440,
     mul_22_8_n_441, mul_22_8_n_442, mul_22_8_n_443, mul_22_8_n_444,
     mul_22_8_n_445, mul_22_8_n_446, mul_22_8_n_447, mul_22_8_n_448,
     mul_22_8_n_449, mul_22_8_n_450, mul_22_8_n_451, mul_22_8_n_452,
     mul_22_8_n_453, mul_22_8_n_454, mul_22_8_n_455, mul_22_8_n_456,
     mul_22_8_n_457, mul_22_8_n_458, mul_22_8_n_459, mul_22_8_n_460,
     mul_22_8_n_461, mul_22_8_n_462, mul_22_8_n_463, mul_22_8_n_464,
     mul_22_8_n_465, mul_22_8_n_466, mul_22_8_n_467, mul_22_8_n_468,
     mul_22_8_n_469, mul_22_8_n_470, mul_22_8_n_471, mul_22_8_n_472,
     mul_22_8_n_473, mul_22_8_n_474, mul_22_8_n_475, mul_22_8_n_476,
     mul_22_8_n_477, mul_22_8_n_478, mul_22_8_n_479, mul_22_8_n_480,
     mul_22_8_n_481, mul_22_8_n_482, mul_22_8_n_483, mul_22_8_n_484,
     mul_22_8_n_485, mul_22_8_n_486, mul_22_8_n_487, mul_22_8_n_488,
     mul_22_8_n_489, mul_22_8_n_490, mul_22_8_n_491, mul_22_8_n_492,
     mul_22_8_n_493, mul_22_8_n_494, mul_22_8_n_495, mul_22_8_n_496,
     mul_22_8_n_497, mul_22_8_n_498, mul_22_8_n_499, mul_22_8_n_500,
     mul_22_8_n_501, mul_22_8_n_502, mul_22_8_n_503, mul_22_8_n_504,
     mul_22_8_n_505, mul_22_8_n_506, mul_22_8_n_507, mul_22_8_n_508,
     mul_22_8_n_509, mul_22_8_n_510, mul_22_8_n_511, mul_22_8_n_512,
     mul_22_8_n_513, mul_22_8_n_514, mul_22_8_n_515, mul_22_8_n_516,
     mul_22_8_n_517, mul_22_8_n_518, mul_22_8_n_519, mul_22_8_n_520,
     mul_22_8_n_521, mul_22_8_n_522, mul_22_8_n_523, mul_22_8_n_524,
     mul_22_8_n_525, mul_22_8_n_526, mul_22_8_n_527, mul_22_8_n_528,
     mul_22_8_n_529, mul_22_8_n_530, mul_22_8_n_531, mul_22_8_n_532,
     mul_22_8_n_533, mul_22_8_n_534, mul_22_8_n_535, mul_22_8_n_536,
     mul_22_8_n_537, mul_22_8_n_538, mul_22_8_n_539, mul_22_8_n_540,
     mul_22_8_n_541, mul_22_8_n_542, mul_22_8_n_543, mul_22_8_n_544,
     mul_22_8_n_545, mul_22_8_n_546, mul_22_8_n_547, mul_22_8_n_548,
     mul_22_8_n_549, mul_22_8_n_550, mul_22_8_n_551, mul_22_8_n_552,
     mul_22_8_n_553, mul_22_8_n_554, mul_22_8_n_555, mul_22_8_n_556,
     mul_22_8_n_557, mul_22_8_n_558, mul_22_8_n_559, mul_22_8_n_560,
     mul_22_8_n_561, mul_22_8_n_562, mul_22_8_n_563, mul_22_8_n_564,
     mul_22_8_n_565, mul_22_8_n_566, mul_22_8_n_567, mul_22_8_n_568,
     mul_22_8_n_569, mul_22_8_n_570, mul_22_8_n_571, mul_22_8_n_572,
     mul_22_8_n_573, mul_22_8_n_574, mul_22_8_n_575, mul_22_8_n_576,
     mul_22_8_n_577, mul_22_8_n_578, mul_22_8_n_579, mul_22_8_n_580,
     mul_22_8_n_581, mul_22_8_n_582, mul_22_8_n_583, mul_22_8_n_584,
     mul_22_8_n_585, mul_22_8_n_586, mul_22_8_n_587, mul_22_8_n_588,
     mul_22_8_n_589, mul_22_8_n_590, mul_22_8_n_591, mul_22_8_n_592,
     mul_22_8_n_593, mul_22_8_n_594, mul_22_8_n_595, mul_22_8_n_596,
     mul_22_8_n_597, mul_22_8_n_598, mul_22_8_n_599, mul_22_8_n_600,
     mul_22_8_n_601, mul_22_8_n_602, mul_22_8_n_603, mul_22_8_n_604,
     mul_22_8_n_605, mul_22_8_n_606, mul_22_8_n_607, mul_22_8_n_608,
     mul_22_8_n_609, mul_22_8_n_610, mul_22_8_n_611, mul_22_8_n_612,
     mul_22_8_n_613, mul_22_8_n_614, mul_22_8_n_615, mul_22_8_n_616,
     mul_22_8_n_617, mul_22_8_n_618, mul_22_8_n_619, mul_22_8_n_620,
     mul_22_8_n_621, mul_22_8_n_622, mul_22_8_n_623, mul_22_8_n_624,
     mul_22_8_n_625, mul_22_8_n_626, mul_22_8_n_627, mul_22_8_n_628,
     mul_22_8_n_629, mul_22_8_n_630, mul_22_8_n_631, mul_22_8_n_632,
     mul_22_8_n_633, mul_22_8_n_634, mul_22_8_n_635, mul_22_8_n_636,
     mul_22_8_n_637, mul_22_8_n_638, mul_22_8_n_639, mul_22_8_n_640,
     mul_22_8_n_641, mul_22_8_n_642, mul_22_8_n_643, mul_22_8_n_644,
     mul_22_8_n_645, mul_22_8_n_646, mul_22_8_n_647, mul_22_8_n_648,
     mul_22_8_n_649, mul_22_8_n_650, mul_22_8_n_651, mul_22_8_n_652,
     mul_22_8_n_653, mul_22_8_n_654, mul_22_8_n_655, mul_22_8_n_656,
     mul_22_8_n_657, mul_22_8_n_658, mul_22_8_n_659, mul_22_8_n_660,
     mul_22_8_n_661, mul_22_8_n_662, mul_22_8_n_663, mul_22_8_n_664,
     mul_22_8_n_665, mul_22_8_n_666, mul_22_8_n_667, mul_22_8_n_668,
     mul_22_8_n_669, mul_22_8_n_670, mul_22_8_n_671, mul_22_8_n_672,
     mul_22_8_n_673, mul_22_8_n_674, mul_22_8_n_675, mul_22_8_n_676,
     mul_22_8_n_677, mul_22_8_n_678, mul_22_8_n_679, mul_22_8_n_680,
     mul_22_8_n_681, mul_22_8_n_682, mul_22_8_n_683, mul_22_8_n_684,
     mul_22_8_n_685, mul_22_8_n_686, mul_22_8_n_688, mul_22_8_n_689,
     mul_22_8_n_690, mul_22_8_n_691, mul_22_8_n_692, mul_22_8_n_693,
     mul_22_8_n_694, mul_22_8_n_695, mul_22_8_n_696, mul_22_8_n_697,
     mul_22_8_n_698, mul_22_8_n_699, mul_22_8_n_700, mul_22_8_n_701,
     mul_22_8_n_702, mul_22_8_n_703, mul_22_8_n_704, mul_22_8_n_705,
     mul_22_8_n_706, mul_22_8_n_707, mul_22_8_n_708, mul_22_8_n_709,
     mul_22_8_n_710, mul_22_8_n_711, mul_22_8_n_712, mul_22_8_n_713,
     mul_22_8_n_714, mul_22_8_n_715, mul_22_8_n_717, mul_22_8_n_718,
     mul_22_8_n_719, mul_22_8_n_720, mul_22_8_n_721, mul_22_8_n_723,
     mul_22_8_n_724, mul_22_8_n_725, mul_22_8_n_726, mul_22_8_n_727,
     mul_22_8_n_728, mul_22_8_n_730, mul_22_8_n_731, mul_22_8_n_732,
     mul_22_8_n_733, mul_22_8_n_734, mul_22_8_n_735, mul_22_8_n_737,
     mul_22_8_n_738, mul_22_8_n_739, mul_22_8_n_740, mul_22_8_n_741,
     mul_22_8_n_742, mul_22_8_n_743, mul_22_8_n_744, mul_22_8_n_745,
     mul_22_8_n_746, mul_22_8_n_747, mul_22_8_n_748, mul_22_8_n_749,
     mul_22_8_n_751, mul_22_8_n_752, mul_22_8_n_754, mul_22_8_n_755,
     mul_22_8_n_756, mul_22_8_n_757, mul_22_8_n_759, mul_22_8_n_760,
     mul_22_8_n_761, mul_22_8_n_762, mul_22_8_n_763, mul_22_8_n_764,
     mul_22_8_n_765, mul_22_8_n_766, mul_22_8_n_767, mul_22_8_n_768,
     mul_22_8_n_769, mul_22_8_n_770, mul_22_8_n_771, mul_22_8_n_772,
     mul_22_8_n_773, mul_22_8_n_774, mul_22_8_n_775, mul_22_8_n_776,
     mul_22_8_n_777, mul_22_8_n_779, mul_22_8_n_780, mul_22_8_n_781,
     mul_22_8_n_782, mul_22_8_n_783, mul_22_8_n_785, mul_22_8_n_786,
     mul_22_8_n_787, mul_22_8_n_788, mul_22_8_n_789, mul_22_8_n_792,
     mul_22_8_n_793, mul_22_8_n_794, mul_22_8_n_795, mul_22_8_n_796,
     mul_22_8_n_797, mul_22_8_n_798, mul_22_8_n_799, mul_22_8_n_800,
     mul_22_8_n_801, mul_22_8_n_802, mul_22_8_n_803, mul_22_8_n_804,
     mul_22_8_n_805, mul_22_8_n_806, mul_22_8_n_807, mul_22_8_n_808,
     mul_22_8_n_809, mul_22_8_n_810, mul_22_8_n_811, mul_22_8_n_812,
     mul_22_8_n_814, mul_22_8_n_815, mul_22_8_n_816, mul_22_8_n_817,
     mul_22_8_n_818, mul_22_8_n_819, mul_22_8_n_821, mul_22_8_n_822,
     mul_22_8_n_823, mul_22_8_n_824, mul_22_8_n_825, mul_22_8_n_826,
     mul_22_8_n_827, mul_22_8_n_828, mul_22_8_n_829, mul_22_8_n_831,
     mul_22_8_n_832, mul_22_8_n_833, mul_22_8_n_834, mul_22_8_n_835,
     mul_22_8_n_836, mul_22_8_n_837, mul_22_8_n_838, mul_22_8_n_839,
     mul_22_8_n_840, mul_22_8_n_841, mul_22_8_n_842, mul_22_8_n_843,
     mul_22_8_n_844, mul_22_8_n_845, mul_22_8_n_846, mul_22_8_n_847,
     mul_22_8_n_848, mul_22_8_n_849, mul_22_8_n_850, mul_22_8_n_851,
     mul_22_8_n_852, mul_22_8_n_853, mul_22_8_n_854, mul_22_8_n_855,
     mul_22_8_n_856, mul_22_8_n_857, mul_22_8_n_858, mul_22_8_n_859,
     mul_22_8_n_860, mul_22_8_n_861, mul_22_8_n_862, mul_22_8_n_863,
     mul_22_8_n_864, mul_22_8_n_867, mul_22_8_n_868, mul_22_8_n_869,
     mul_22_8_n_870, mul_22_8_n_871, mul_22_8_n_872, mul_22_8_n_873,
     mul_22_8_n_874, mul_22_8_n_875, mul_22_8_n_877, mul_22_8_n_879,
     mul_22_8_n_880, mul_22_8_n_881, mul_22_8_n_882, mul_22_8_n_883,
     mul_22_8_n_884, mul_22_8_n_885, mul_22_8_n_886, mul_22_8_n_887,
     mul_22_8_n_888, mul_22_8_n_889, mul_22_8_n_892, mul_22_8_n_893,
     mul_22_8_n_894, mul_22_8_n_895, mul_22_8_n_897, mul_22_8_n_898,
     mul_22_8_n_903, mul_22_8_n_904, mul_22_8_n_908, mul_22_8_n_911,
     mul_22_8_n_912, mul_22_8_n_913, mul_22_8_n_914, mul_22_8_n_915,
     mul_22_8_n_916, mul_22_8_n_917, mul_22_8_n_918, mul_22_8_n_919,
     mul_22_8_n_920, mul_22_8_n_921, mul_22_8_n_922, mul_22_8_n_923,
     mul_22_8_n_924, mul_22_8_n_925, mul_22_8_n_926, mul_22_8_n_927,
     mul_22_8_n_928, mul_22_8_n_929, mul_22_8_n_930, mul_22_8_n_931,
     mul_22_8_n_932, mul_22_8_n_933, mul_22_8_n_934, mul_22_8_n_935,
     mul_22_8_n_936, mul_22_8_n_937, mul_22_8_n_938, mul_22_8_n_939,
     mul_22_8_n_940, mul_22_8_n_941, mul_22_8_n_942, mul_22_8_n_943,
     mul_22_8_n_944, mul_22_8_n_945, mul_22_8_n_946, mul_22_8_n_947,
     mul_22_8_n_948, mul_22_8_n_949, mul_22_8_n_950, mul_22_8_n_951,
     mul_22_8_n_952, mul_22_8_n_953, mul_22_8_n_954, mul_22_8_n_955,
     mul_22_8_n_956, mul_22_8_n_957, mul_22_8_n_958, mul_22_8_n_959,
     mul_22_8_n_960, mul_22_8_n_961, mul_22_8_n_962, mul_22_8_n_963,
     mul_22_8_n_964, mul_22_8_n_965, mul_22_8_n_966, mul_22_8_n_967,
     mul_22_8_n_968, mul_22_8_n_969, mul_22_8_n_970, mul_22_8_n_971,
     mul_22_8_n_972, mul_22_8_n_973, mul_22_8_n_974, mul_22_8_n_975,
     mul_22_8_n_976, mul_22_8_n_977, mul_22_8_n_978, mul_22_8_n_979,
     mul_22_8_n_980, mul_22_8_n_981, mul_22_8_n_982, mul_22_8_n_983,
     mul_22_8_n_984, mul_22_8_n_985, mul_22_8_n_986, mul_22_8_n_987,
     mul_22_8_n_988, mul_22_8_n_989, mul_22_8_n_990, mul_22_8_n_991,
     mul_22_8_n_992, mul_22_8_n_993, mul_22_8_n_994, mul_22_8_n_995,
     mul_22_8_n_996, mul_22_8_n_997, mul_22_8_n_998, mul_22_8_n_999,
     mul_22_8_n_1000, mul_22_8_n_1001, mul_22_8_n_1002, mul_22_8_n_1003,
     mul_22_8_n_1004, mul_22_8_n_1005, mul_22_8_n_1006, mul_22_8_n_1007,
     mul_22_8_n_1008, mul_22_8_n_1009, mul_22_8_n_1010, mul_22_8_n_1011,
     mul_22_8_n_1012, mul_22_8_n_1013, mul_22_8_n_1014, mul_22_8_n_1015,
     mul_22_8_n_1016, mul_22_8_n_1017, mul_22_8_n_1018, mul_22_8_n_1019,
     mul_22_8_n_1020, mul_22_8_n_1021, mul_22_8_n_1022, mul_22_8_n_1023,
     mul_22_8_n_1024, mul_22_8_n_1025, mul_22_8_n_1026, mul_22_8_n_1027,
     mul_22_8_n_1028, mul_22_8_n_1029, mul_22_8_n_1030, mul_22_8_n_1031,
     mul_22_8_n_1032, mul_22_8_n_1033, mul_22_8_n_1034, mul_22_8_n_1035,
     mul_22_8_n_1036, mul_22_8_n_1037, mul_22_8_n_1038, mul_22_8_n_1039,
     mul_22_8_n_1040, mul_22_8_n_1041, mul_22_8_n_1042, mul_22_8_n_1043,
     mul_22_8_n_1044, mul_22_8_n_1045, mul_22_8_n_1046, mul_22_8_n_1047,
     mul_22_8_n_1048, mul_22_8_n_1049, mul_22_8_n_1050, mul_22_8_n_1051,
     mul_22_8_n_1052, mul_22_8_n_1053, mul_22_8_n_1054, mul_22_8_n_1055,
     mul_22_8_n_1056, mul_22_8_n_1057, mul_22_8_n_1058, mul_22_8_n_1059,
     mul_22_8_n_1060, mul_22_8_n_1061, mul_22_8_n_1062, mul_22_8_n_1063,
     mul_22_8_n_1064, mul_22_8_n_1065, mul_22_8_n_1066, mul_22_8_n_1067,
     mul_22_8_n_1068, mul_22_8_n_1069, mul_22_8_n_1070, mul_22_8_n_1071,
     mul_22_8_n_1072, mul_22_8_n_1073, mul_22_8_n_1074, mul_22_8_n_1075,
     mul_22_8_n_1076, mul_22_8_n_1077, mul_22_8_n_1078, mul_22_8_n_1079,
     mul_22_8_n_1080, mul_22_8_n_1081, mul_22_8_n_1082, mul_22_8_n_1083,
     mul_22_8_n_1084, mul_22_8_n_1085, mul_22_8_n_1086, mul_22_8_n_1087,
     mul_22_8_n_1088, mul_22_8_n_1089, mul_22_8_n_1090, mul_22_8_n_1091,
     mul_22_8_n_1092, mul_22_8_n_1093, mul_22_8_n_1094, mul_22_8_n_1095,
     mul_22_8_n_1096, mul_22_8_n_1097, mul_22_8_n_1098, mul_22_8_n_1099,
     mul_22_8_n_1100, mul_22_8_n_1101, mul_22_8_n_1102, mul_22_8_n_1103,
     mul_22_8_n_1104, mul_22_8_n_1105, mul_22_8_n_1106, mul_22_8_n_1107,
     mul_22_8_n_1108, mul_22_8_n_1109, mul_22_8_n_1110, mul_22_8_n_1111,
     mul_22_8_n_1112, mul_22_8_n_1113, mul_22_8_n_1114, mul_22_8_n_1115,
     mul_22_8_n_1116, mul_22_8_n_1117, mul_22_8_n_1118, mul_22_8_n_1119,
     mul_22_8_n_1120, mul_22_8_n_1121, mul_22_8_n_1122, mul_22_8_n_1123,
     mul_22_8_n_1124, mul_22_8_n_1125, mul_22_8_n_1126, mul_22_8_n_1127,
     mul_22_8_n_1128, mul_22_8_n_1129, mul_22_8_n_1130, mul_22_8_n_1131,
     mul_22_8_n_1132, mul_22_8_n_1133, mul_22_8_n_1134, mul_22_8_n_1135,
     mul_22_8_n_1136, mul_22_8_n_1137, mul_22_8_n_1138, mul_22_8_n_1139,
     mul_22_8_n_1140, mul_22_8_n_1141, mul_22_8_n_1142, mul_22_8_n_1143,
     mul_22_8_n_1144, mul_22_8_n_1145, mul_22_8_n_1146, mul_22_8_n_1147,
     mul_22_8_n_1148, mul_22_8_n_1149, mul_22_8_n_1150, mul_22_8_n_1151,
     mul_22_8_n_1152, mul_22_8_n_1153, mul_22_8_n_1154, mul_22_8_n_1155,
     mul_22_8_n_1156, mul_22_8_n_1157, mul_22_8_n_1158, mul_22_8_n_1159,
     mul_22_8_n_1160, mul_22_8_n_1161, mul_22_8_n_1162, mul_22_8_n_1163,
     mul_22_8_n_1164, mul_22_8_n_1165, mul_22_8_n_1166, mul_22_8_n_1167,
     mul_22_8_n_1168, mul_22_8_n_1169, mul_22_8_n_1170, mul_22_8_n_1171,
     mul_22_8_n_1172, mul_22_8_n_1173, mul_22_8_n_1174, mul_22_8_n_1175,
     mul_22_8_n_1176, mul_22_8_n_1177, mul_22_8_n_1178, mul_22_8_n_1179,
     mul_22_8_n_1180, mul_22_8_n_1181, mul_22_8_n_1182, mul_22_8_n_1183,
     mul_22_8_n_1184, mul_22_8_n_1185, mul_22_8_n_1186, mul_22_8_n_1187,
     mul_22_8_n_1188, mul_22_8_n_1189, mul_22_8_n_1190, mul_22_8_n_1191,
     mul_22_8_n_1192, mul_22_8_n_1193, mul_22_8_n_1194, mul_22_8_n_1195,
     mul_22_8_n_1196, mul_22_8_n_1197, mul_22_8_n_1198, mul_22_8_n_1199,
     mul_22_8_n_1200, mul_22_8_n_1201, mul_22_8_n_1202, mul_22_8_n_1203,
     mul_22_8_n_1204, mul_22_8_n_1205, mul_22_8_n_1206, mul_22_8_n_1207,
     mul_22_8_n_1208, mul_22_8_n_1209, mul_22_8_n_1210, mul_22_8_n_1211,
     mul_22_8_n_1212, mul_22_8_n_1213, mul_22_8_n_1214, mul_22_8_n_1215,
     mul_22_8_n_1216, mul_22_8_n_1217, mul_22_8_n_1218, mul_22_8_n_1219,
     mul_22_8_n_1220, mul_22_8_n_1221, mul_22_8_n_1222, mul_22_8_n_1223,
     mul_22_8_n_1224, mul_22_8_n_1225, mul_22_8_n_1226, mul_22_8_n_1227,
     mul_22_8_n_1228, mul_22_8_n_1229, mul_22_8_n_1230, mul_22_8_n_1231,
     mul_22_8_n_1232, mul_22_8_n_1233, mul_22_8_n_1234, mul_22_8_n_1235,
     mul_22_8_n_1236, mul_22_8_n_1237, mul_22_8_n_1238, mul_22_8_n_1239,
     mul_22_8_n_1240, mul_22_8_n_1241, mul_22_8_n_1242, mul_22_8_n_1243,
     mul_22_8_n_1244, mul_22_8_n_1245, mul_22_8_n_1246, mul_22_8_n_1247,
     mul_22_8_n_1248, mul_22_8_n_1249, mul_22_8_n_1250, mul_22_8_n_1251,
     mul_22_8_n_1252, mul_22_8_n_1253, mul_22_8_n_1254, mul_22_8_n_1255,
     mul_22_8_n_1256, mul_22_8_n_1257, mul_22_8_n_1258, mul_22_8_n_1259,
     mul_22_8_n_1260, mul_22_8_n_1261, mul_22_8_n_1262, mul_22_8_n_1263,
     mul_22_8_n_1264, mul_22_8_n_1265, mul_22_8_n_1266, mul_22_8_n_1267,
     mul_22_8_n_1268, mul_22_8_n_1269, mul_22_8_n_1270, mul_22_8_n_1271,
     mul_22_8_n_1272, mul_22_8_n_1273, mul_22_8_n_1274, mul_22_8_n_1275,
     mul_22_8_n_1276, mul_22_8_n_1277, mul_22_8_n_1278, mul_22_8_n_1279,
     mul_22_8_n_1280, mul_22_8_n_1281, mul_22_8_n_1282, mul_22_8_n_1283,
     mul_22_8_n_1284, mul_22_8_n_1285, mul_22_8_n_1286, mul_22_8_n_1287,
     mul_22_8_n_1288, mul_22_8_n_1289, mul_22_8_n_1290, mul_22_8_n_1291,
     mul_22_8_n_1292, mul_22_8_n_1293, mul_22_8_n_1294, mul_22_8_n_1295,
     mul_22_8_n_1296, mul_22_8_n_1297, mul_22_8_n_1298, mul_22_8_n_1299,
     mul_22_8_n_1300, mul_22_8_n_1301, mul_22_8_n_1302, mul_22_8_n_1303,
     mul_22_8_n_1304, mul_22_8_n_1305, mul_22_8_n_1306, mul_22_8_n_1307,
     mul_22_8_n_1308, mul_22_8_n_1309, mul_22_8_n_1310, mul_22_8_n_1311,
     mul_22_8_n_1312, mul_22_8_n_1313, mul_22_8_n_1314, mul_22_8_n_1315,
     mul_22_8_n_1316, n_0, n_23, n_24, n_25, n_26, n_27, n_28, n_31, n_34, n_35,
     n_36, n_37, n_38, n_40, n_42, n_43, n_44, n_45, n_46, n_47, n_48, n_49,
     n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58, n_59, n_60, n_61,
     n_62, n_63, n_64, n_65, n_66, n_67, n_68, n_69, n_70, n_72, n_73, n_74,
     n_75, n_77, n_78, n_80, n_81, n_84, n_85, n_86, clk, clr, n_154, n_155,
     asc001_0_, asc001_1_, asc001_2_, asc001_3_, asc001_4_, asc001_5_, asc001_6_,
     asc001_7_, asc001_8_, asc001_9_, asc001_10_, asc001_11_, asc001_12_,
     asc001_13_, asc001_14_, asc001_15_, asc001_16_, asc001_17_, asc001_18_,
     asc001_19_, asc001_20_, asc001_21_, asc001_22_, asc001_23_, asc001_24_,
     asc001_25_, asc001_26_, asc001_27_, asc001_28_, asc001_29_, asc001_30_,
     asc001_31_;
assign {out1[31]} = asc001_31_;
assign {out1[30]} = asc001_30_;
assign {out1[29]} = asc001_29_;
assign {out1[28]} = asc001_28_;
assign {out1[27]} = asc001_27_;
assign {out1[26]} = asc001_26_;
assign {out1[25]} = asc001_25_;
assign {out1[24]} = asc001_24_;
assign {out1[23]} = asc001_23_;
assign {out1[22]} = asc001_22_;
assign {out1[21]} = asc001_21_;
assign {out1[20]} = asc001_20_;
assign {out1[19]} = asc001_19_;
assign {out1[18]} = asc001_18_;
assign {out1[17]} = asc001_17_;
assign {out1[16]} = asc001_16_;
assign {out1[15]} = asc001_15_;
assign {out1[14]} = asc001_14_;
assign {out1[13]} = asc001_13_;
assign {out1[12]} = asc001_12_;
assign {out1[11]} = asc001_11_;
assign {out1[10]} = asc001_10_;
 reg retime_s1_13_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_13_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_13_reg_reg_IQ <= mul_22_8_n_1283;
     end
 assign n_72 = retime_s1_13_reg_reg_IQ;
 reg out1_23_L0_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) out1_23_L0_reg_IQ <= 1'B0;
     else begin
         out1_23_L0_reg_IQ <= asc001_8_;
     end
 assign {out1[8]} = out1_23_L0_reg_IQ;
 reg out1_24_L0_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) out1_24_L0_reg_IQ <= 1'B0;
     else begin
         out1_24_L0_reg_IQ <= asc001_7_;
     end
 assign {out1[7]} = out1_24_L0_reg_IQ;
 reg out1_25_L0_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) out1_25_L0_reg_IQ <= 1'B0;
     else begin
         out1_25_L0_reg_IQ <= asc001_6_;
     end
 assign {out1[6]} = out1_25_L0_reg_IQ;
 reg out1_26_L0_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) out1_26_L0_reg_IQ <= 1'B0;
     else begin
         out1_26_L0_reg_IQ <= asc001_5_;
     end
 assign {out1[5]} = out1_26_L0_reg_IQ;
 reg out1_27_L0_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) out1_27_L0_reg_IQ <= 1'B0;
     else begin
         out1_27_L0_reg_IQ <= asc001_4_;
     end
 assign {out1[4]} = out1_27_L0_reg_IQ;
 reg out1_28_L0_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) out1_28_L0_reg_IQ <= 1'B0;
     else begin
         out1_28_L0_reg_IQ <= asc001_3_;
     end
 assign {out1[3]} = out1_28_L0_reg_IQ;
 reg out1_29_L0_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) out1_29_L0_reg_IQ <= 1'B0;
     else begin
         out1_29_L0_reg_IQ <= asc001_2_;
     end
 assign {out1[2]} = out1_29_L0_reg_IQ;
 reg out1_30_L0_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) out1_30_L0_reg_IQ <= 1'B0;
     else begin
         out1_30_L0_reg_IQ <= asc001_1_;
     end
 assign {out1[1]} = out1_30_L0_reg_IQ;
 reg out1_31_L0_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) out1_31_L0_reg_IQ <= 1'B0;
     else begin
         out1_31_L0_reg_IQ <= asc001_0_;
     end
 assign {out1[0]} = out1_31_L0_reg_IQ;
 reg retime_s1_1_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_1_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_1_reg_reg_IQ <= mul_22_8_n_779;
     end
 assign n_86 = retime_s1_1_reg_reg_IQ;
 reg retime_s1_7_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_7_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_7_reg_reg_IQ <= mul_22_8_n_825;
     end
 assign n_78 = retime_s1_7_reg_reg_IQ;
 reg retime_s1_10_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_10_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_10_reg_reg_IQ <= mul_22_8_n_822;
     end
 assign n_75 = retime_s1_10_reg_reg_IQ;
 reg retime_s1_11_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_11_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_11_reg_reg_IQ <= mul_22_8_n_1100;
     end
 assign n_74 = retime_s1_11_reg_reg_IQ;
 reg out1_22_L0_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) out1_22_L0_reg_IQ <= 1'B0;
     else begin
         out1_22_L0_reg_IQ <= asc001_9_;
     end
 assign {out1[9]} = out1_22_L0_reg_IQ;
 reg retime_s1_15_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_15_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_15_reg_reg_IQ <= mul_22_8_n_1018;
     end
 assign n_69 = retime_s1_15_reg_reg_IQ;
 reg retime_s1_20_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_20_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_20_reg_reg_IQ <= mul_22_8_n_769;
     end
 assign n_64 = retime_s1_20_reg_reg_IQ;
 reg retime_s1_27_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_27_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_27_reg_reg_IQ <= mul_22_8_n_1135;
     end
 assign n_57 = retime_s1_27_reg_reg_IQ;
 reg retime_s1_28_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_28_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_28_reg_reg_IQ <= mul_22_8_n_971;
     end
 assign n_56 = retime_s1_28_reg_reg_IQ;
 reg retime_s1_30_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_30_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_30_reg_reg_IQ <= mul_22_8_n_945;
     end
 assign n_54 = retime_s1_30_reg_reg_IQ;
 reg retime_s1_33_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_33_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_33_reg_reg_IQ <= mul_22_8_n_920;
     end
 assign n_51 = retime_s1_33_reg_reg_IQ;
 reg retime_s1_36_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_36_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_36_reg_reg_IQ <= mul_22_8_n_815;
     end
 assign n_48 = retime_s1_36_reg_reg_IQ;
 reg retime_s1_37_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_37_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_37_reg_reg_IQ <= mul_22_8_n_794;
     end
 assign n_47 = retime_s1_37_reg_reg_IQ;
 reg retime_s1_38_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_38_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_38_reg_reg_IQ <= mul_22_8_n_797;
     end
 assign n_46 = retime_s1_38_reg_reg_IQ;
 reg retime_s1_40_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_40_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_40_reg_reg_IQ <= mul_22_8_n_995;
     end
 assign n_44 = retime_s1_40_reg_reg_IQ;
 reg retime_s1_43_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_43_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_43_reg_reg_IQ <= mul_22_8_n_1061;
     end
 assign n_40 = retime_s1_43_reg_reg_IQ;
 reg retime_s1_44_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_44_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_44_reg_reg_IQ <= mul_22_8_n_2;
     end
 assign n_38 = retime_s1_44_reg_reg_IQ;
 reg retime_s1_46_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_46_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_46_reg_reg_IQ <= mul_22_8_n_1281;
     end
 assign n_36 = retime_s1_46_reg_reg_IQ;
 reg retime_s1_48_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_48_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_48_reg_reg_IQ <= mul_22_8_n_781;
     end
 assign n_34 = retime_s1_48_reg_reg_IQ;
 reg retime_s1_49_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_49_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_49_reg_reg_IQ <= mul_22_8_n_798;
     end
 assign n_31 = retime_s1_49_reg_reg_IQ;
 reg retime_s1_21_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_21_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_21_reg_reg_IQ <= mul_22_8_n_780;
     end
 assign n_63 = retime_s1_21_reg_reg_IQ;
 reg retime_s1_51_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_51_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_51_reg_reg_IQ <= mul_22_8_n_777;
     end
 assign n_27 = retime_s1_51_reg_reg_IQ;
 reg retime_s1_52_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_52_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_52_reg_reg_IQ <= mul_22_8_n_796;
     end
 assign n_26 = retime_s1_52_reg_reg_IQ;
 reg retime_s1_39_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_39_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_39_reg_reg_IQ <= mul_22_8_n_799;
     end
 assign n_45 = retime_s1_39_reg_reg_IQ;
 reg retime_s1_3_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_3_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_3_reg_reg_IQ <= mul_22_8_n_996;
     end
 assign n_84 = retime_s1_3_reg_reg_IQ;
 reg retime_s1_4_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_4_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_4_reg_reg_IQ <= mul_22_8_n_1305;
     end
 assign n_81 = retime_s1_4_reg_reg_IQ;
 reg retime_s1_47_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_47_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_47_reg_reg_IQ <= mul_22_8_n_1136;
     end
 assign n_35 = retime_s1_47_reg_reg_IQ;
 reg retime_s1_5_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_5_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_5_reg_reg_IQ <= mul_22_8_n_1099;
     end
 assign n_80 = retime_s1_5_reg_reg_IQ;
 reg retime_s1_2_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_2_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_2_reg_reg_IQ <= mul_22_8_n_972;
     end
 assign n_85 = retime_s1_2_reg_reg_IQ;
 reg retime_s1_8_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_8_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_8_reg_reg_IQ <= mul_22_8_n_1134;
     end
 assign n_77 = retime_s1_8_reg_reg_IQ;
 reg retime_s1_12_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_12_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_12_reg_reg_IQ <= mul_22_8_n_1308;
     end
 assign n_73 = retime_s1_12_reg_reg_IQ;
 reg retime_s1_14_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_14_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_14_reg_reg_IQ <= mul_22_8_n_1062;
     end
 assign n_70 = retime_s1_14_reg_reg_IQ;
 reg retime_s1_42_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_42_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_42_reg_reg_IQ <= mul_22_8_n_792;
     end
 assign n_42 = retime_s1_42_reg_reg_IQ;
 reg retime_s1_16_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_16_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_16_reg_reg_IQ <= mul_22_8_n_921;
     end
 assign n_68 = retime_s1_16_reg_reg_IQ;
 reg retime_s1_18_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_18_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_18_reg_reg_IQ <= mul_22_8_n_782;
     end
 assign n_66 = retime_s1_18_reg_reg_IQ;
 reg retime_s1_19_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_19_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_19_reg_reg_IQ <= mul_22_8_n_766;
     end
 assign n_65 = retime_s1_19_reg_reg_IQ;
 reg retime_s1_50_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_50_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_50_reg_reg_IQ <= mul_22_8_n_831;
     end
 assign n_28 = retime_s1_50_reg_reg_IQ;
 reg retime_s1_22_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_22_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_22_reg_reg_IQ <= mul_22_8_n_795;
     end
 assign n_62 = retime_s1_22_reg_reg_IQ;
 reg retime_s1_23_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_23_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_23_reg_reg_IQ <= mul_22_8_n_801;
     end
 assign n_61 = retime_s1_23_reg_reg_IQ;
 reg retime_s1_17_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_17_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_17_reg_reg_IQ <= mul_22_8_n_763;
     end
 assign n_67 = retime_s1_17_reg_reg_IQ;
 reg retime_s1_25_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_25_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_25_reg_reg_IQ <= mul_22_8_n_1060;
     end
 assign n_59 = retime_s1_25_reg_reg_IQ;
 reg retime_s1_26_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_26_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_26_reg_reg_IQ <= mul_22_8_n_1101;
     end
 assign n_58 = retime_s1_26_reg_reg_IQ;
 reg retime_s1_29_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_29_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_29_reg_reg_IQ <= mul_22_8_n_994;
     end
 assign n_55 = retime_s1_29_reg_reg_IQ;
 reg retime_s1_31_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_31_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_31_reg_reg_IQ <= mul_22_8_n_970;
     end
 assign n_53 = retime_s1_31_reg_reg_IQ;
 reg retime_s1_34_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_34_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_34_reg_reg_IQ <= mul_22_8_n_793;
     end
 assign n_50 = retime_s1_34_reg_reg_IQ;
 reg retime_s1_35_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_35_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_35_reg_reg_IQ <= mul_22_8_n_816;
     end
 assign n_49 = retime_s1_35_reg_reg_IQ;
 reg retime_s1_32_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_32_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_32_reg_reg_IQ <= mul_22_8_n_947;
     end
 assign n_52 = retime_s1_32_reg_reg_IQ;
 reg retime_s1_41_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_41_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_41_reg_reg_IQ <= mul_22_8_n_1017;
     end
 assign n_43 = retime_s1_41_reg_reg_IQ;
 reg retime_s1_45_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_45_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_45_reg_reg_IQ <= mul_22_8_n_1306;
     end
 assign n_37 = retime_s1_45_reg_reg_IQ;
 reg retime_s1_24_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_24_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_24_reg_reg_IQ <= mul_22_8_n_800;
     end
 assign n_60 = retime_s1_24_reg_reg_IQ;
 reg retime_s1_53_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_53_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_53_reg_reg_IQ <= mul_22_8_n_919;
     end
 assign n_25 = retime_s1_53_reg_reg_IQ;
 reg retime_s1_54_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_54_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_54_reg_reg_IQ <= mul_22_8_n_946;
     end
 assign n_24 = retime_s1_54_reg_reg_IQ;
 reg retime_s1_55_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_55_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_55_reg_reg_IQ <= mul_22_8_n_1019;
     end
 assign n_23 = retime_s1_55_reg_reg_IQ;
 reg retime_s1_9_reg_reg_IQ;
 wire retime_s1_9_reg_reg_IQN;
 assign retime_s1_9_reg_reg_IQN = !retime_s1_9_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_9_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_9_reg_reg_IQ <= mul_22_8_n_1287;
     end
 assign mul_22_8_n_828 = retime_s1_9_reg_reg_IQN;
 reg retime_s1_6_reg_reg_IQ;
 wire retime_s1_6_reg_reg_IQN;
 assign retime_s1_6_reg_reg_IQN = !retime_s1_6_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_6_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_6_reg_reg_IQ <= mul_22_8_n_1285;
     end
 assign mul_22_8_n_823 = retime_s1_6_reg_reg_IQN;
 assign mul_22_8_n_918 = ((mul_22_8_n_477 & mul_22_8_n_391) | (mul_22_8_n_421 & (mul_22_8_n_477 ^ mul_22_8_n_391)));
 assign mul_22_8_n_917 = (mul_22_8_n_421 ^ (mul_22_8_n_477 ^ mul_22_8_n_391));
 assign mul_22_8_n_1293 = ((mul_22_8_n_618 & mul_22_8_n_519) | (mul_22_8_n_706 & (mul_22_8_n_618 ^ mul_22_8_n_519)));
 assign mul_22_8_n_916 = (mul_22_8_n_706 ^ (mul_22_8_n_618 ^ mul_22_8_n_519));
 assign mul_22_8_n_1268 = ((mul_22_8_n_397 & mul_22_8_n_385) | (mul_22_8_n_513 & (mul_22_8_n_397 ^ mul_22_8_n_385)));
 assign mul_22_8_n_1269 = (mul_22_8_n_513 ^ (mul_22_8_n_397 ^ mul_22_8_n_385));
 assign mul_22_8_n_915 = ((mul_22_8_n_692 & mul_22_8_n_557) | (mul_22_8_n_1269 & (mul_22_8_n_692 ^ mul_22_8_n_557)));
 assign mul_22_8_n_914 = (mul_22_8_n_1269 ^ (mul_22_8_n_692 ^ mul_22_8_n_557));
 assign mul_22_8_n_1266 = ((mul_22_8_n_566 & mul_22_8_n_620) | (mul_22_8_n_582 & (mul_22_8_n_566 ^ mul_22_8_n_620)));
 assign mul_22_8_n_1267 = (mul_22_8_n_582 ^ (mul_22_8_n_566 ^ mul_22_8_n_620));
 assign mul_22_8_n_913 = ((mul_22_8_n_1268 & mul_22_8_n_704) | (mul_22_8_n_1267 & (mul_22_8_n_1268 ^
    mul_22_8_n_704)));
 assign mul_22_8_n_912 = (mul_22_8_n_1267 ^ (mul_22_8_n_1268 ^ mul_22_8_n_704));
 assign mul_22_8_n_1263 = ((mul_22_8_n_400 & mul_22_8_n_384) | (mul_22_8_n_551 & (mul_22_8_n_400 ^ mul_22_8_n_384)));
 assign mul_22_8_n_1265 = (mul_22_8_n_551 ^ (mul_22_8_n_400 ^ mul_22_8_n_384));
 assign mul_22_8_n_1261 = ((mul_22_8_n_541 & mul_22_8_n_542) | (mul_22_8_n_694 & (mul_22_8_n_541 ^ mul_22_8_n_542)));
 assign mul_22_8_n_1264 = (mul_22_8_n_694 ^ (mul_22_8_n_541 ^ mul_22_8_n_542));
 assign mul_22_8_n_1294 = ((mul_22_8_n_1265 & mul_22_8_n_1266) | (mul_22_8_n_1264 & (mul_22_8_n_1265
    ^ mul_22_8_n_1266)));
 assign mul_22_8_n_911 = (mul_22_8_n_1264 ^ (mul_22_8_n_1265 ^ mul_22_8_n_1266));
 assign mul_22_8_n_1259 = ((mul_22_8_n_621 & mul_22_8_n_619) | (mul_22_8_n_410 & (mul_22_8_n_621 ^ mul_22_8_n_619)));
 assign mul_22_8_n_1262 = (mul_22_8_n_410 ^ (mul_22_8_n_621 ^ mul_22_8_n_619));
 assign mul_22_8_n_1256 = ((mul_22_8_n_711 & mul_22_8_n_510) | (mul_22_8_n_1263 & (mul_22_8_n_711 ^ mul_22_8_n_510)));
 assign mul_22_8_n_1260 = (mul_22_8_n_1263 ^ (mul_22_8_n_711 ^ mul_22_8_n_510));
 assign mul_22_8_n_1295 = ((mul_22_8_n_1261 & mul_22_8_n_1262) | (mul_22_8_n_1260 & (mul_22_8_n_1261
    ^ mul_22_8_n_1262)));
 assign mul_22_8_n_1270 = (mul_22_8_n_1260 ^ (mul_22_8_n_1261 ^ mul_22_8_n_1262));
 assign mul_22_8_n_1254 = ((mul_22_8_n_492 & mul_22_8_n_388) | (mul_22_8_n_490 & (mul_22_8_n_492 ^ mul_22_8_n_388)));
 assign mul_22_8_n_1258 = (mul_22_8_n_490 ^ (mul_22_8_n_492 ^ mul_22_8_n_388));
 assign mul_22_8_n_1253 = ((mul_22_8_n_402 & mul_22_8_n_539) | (mul_22_8_n_571 & (mul_22_8_n_402 ^ mul_22_8_n_539)));
 assign mul_22_8_n_1257 = (mul_22_8_n_571 ^ (mul_22_8_n_402 ^ mul_22_8_n_539));
 assign mul_22_8_n_1249 = ((mul_22_8_n_1259 & mul_22_8_n_686) | (mul_22_8_n_1258 & (mul_22_8_n_1259 ^
    mul_22_8_n_686)));
 assign mul_22_8_n_1255 = (mul_22_8_n_1258 ^ (mul_22_8_n_1259 ^ mul_22_8_n_686));
 assign mul_22_8_n_1296 = ((mul_22_8_n_1256 & mul_22_8_n_1257) | (mul_22_8_n_1255 & (mul_22_8_n_1256
    ^ mul_22_8_n_1257)));
 assign mul_22_8_n_1271 = (mul_22_8_n_1255 ^ (mul_22_8_n_1256 ^ mul_22_8_n_1257));
 assign mul_22_8_n_1248 = ((mul_22_8_n_458 & mul_22_8_n_462) | (mul_22_8_n_401 & (mul_22_8_n_458 ^ mul_22_8_n_462)));
 assign mul_22_8_n_1252 = (mul_22_8_n_401 ^ (mul_22_8_n_458 ^ mul_22_8_n_462));
 assign mul_22_8_n_1245 = ((mul_22_8_n_494 & mul_22_8_n_622) | (mul_22_8_n_709 & (mul_22_8_n_494 ^ mul_22_8_n_622)));
 assign mul_22_8_n_1251 = (mul_22_8_n_709 ^ (mul_22_8_n_494 ^ mul_22_8_n_622));
 assign mul_22_8_n_1243 = ((mul_22_8_n_1253 & mul_22_8_n_1254) | (mul_22_8_n_1252 & (mul_22_8_n_1253
    ^ mul_22_8_n_1254)));
 assign mul_22_8_n_1250 = (mul_22_8_n_1252 ^ (mul_22_8_n_1253 ^ mul_22_8_n_1254));
 assign mul_22_8_n_1297 = ((mul_22_8_n_1250 & mul_22_8_n_1251) | (mul_22_8_n_1249 & (mul_22_8_n_1250
    ^ mul_22_8_n_1251)));
 assign mul_22_8_n_1272 = (mul_22_8_n_1249 ^ (mul_22_8_n_1250 ^ mul_22_8_n_1251));
 assign mul_22_8_n_1241 = ((mul_22_8_n_616 & mul_22_8_n_386) | (mul_22_8_n_611 & (mul_22_8_n_616 ^ mul_22_8_n_386)));
 assign mul_22_8_n_1246 = (mul_22_8_n_611 ^ (mul_22_8_n_616 ^ mul_22_8_n_386));
 assign mul_22_8_n_1240 = ((mul_22_8_n_405 & mul_22_8_n_605) | (mul_22_8_n_599 & (mul_22_8_n_405 ^ mul_22_8_n_605)));
 assign mul_22_8_n_1247 = (mul_22_8_n_599 ^ (mul_22_8_n_405 ^ mul_22_8_n_605));
 assign mul_22_8_n_1237 = ((mul_22_8_n_685 & mul_22_8_n_576) | (mul_22_8_n_1248 & (mul_22_8_n_685 ^ mul_22_8_n_576)));
 assign mul_22_8_n_1244 = (mul_22_8_n_1248 ^ (mul_22_8_n_685 ^ mul_22_8_n_576));
 assign mul_22_8_n_1235 = ((mul_22_8_n_1246 & mul_22_8_n_1247) | (mul_22_8_n_1245 & (mul_22_8_n_1246
    ^ mul_22_8_n_1247)));
 assign mul_22_8_n_1242 = (mul_22_8_n_1245 ^ (mul_22_8_n_1246 ^ mul_22_8_n_1247));
 assign mul_22_8_n_1298 = ((mul_22_8_n_1243 & mul_22_8_n_1244) | (mul_22_8_n_1242 & (mul_22_8_n_1243
    ^ mul_22_8_n_1244)));
 assign mul_22_8_n_1273 = (mul_22_8_n_1242 ^ (mul_22_8_n_1243 ^ mul_22_8_n_1244));
 assign mul_22_8_n_1233 = ((mul_22_8_n_590 & mul_22_8_n_651) | (mul_22_8_n_534 & (mul_22_8_n_590 ^ mul_22_8_n_651)));
 assign mul_22_8_n_1238 = (mul_22_8_n_534 ^ (mul_22_8_n_590 ^ mul_22_8_n_651));
 assign mul_22_8_n_1232 = ((mul_22_8_n_567 & mul_22_8_n_658) | (mul_22_8_n_623 & (mul_22_8_n_567 ^ mul_22_8_n_658)));
 assign mul_22_8_n_1239 = (mul_22_8_n_623 ^ (mul_22_8_n_567 ^ mul_22_8_n_658));
 assign mul_22_8_n_1228 = ((mul_22_8_n_1241 & mul_22_8_n_703) | (mul_22_8_n_1240 & (mul_22_8_n_1241 ^
    mul_22_8_n_703)));
 assign mul_22_8_n_1236 = (mul_22_8_n_1240 ^ (mul_22_8_n_1241 ^ mul_22_8_n_703));
 assign mul_22_8_n_1225 = ((mul_22_8_n_1238 & mul_22_8_n_1239) | (mul_22_8_n_1237 & (mul_22_8_n_1238
    ^ mul_22_8_n_1239)));
 assign mul_22_8_n_1234 = (mul_22_8_n_1237 ^ (mul_22_8_n_1238 ^ mul_22_8_n_1239));
 assign mul_22_8_n_1299 = ((mul_22_8_n_1235 & mul_22_8_n_1236) | (mul_22_8_n_1234 & (mul_22_8_n_1235
    ^ mul_22_8_n_1236)));
 assign mul_22_8_n_1274 = (mul_22_8_n_1234 ^ (mul_22_8_n_1235 ^ mul_22_8_n_1236));
 assign mul_22_8_n_1224 = ((mul_22_8_n_396 & mul_22_8_n_387) | (mul_22_8_n_653 & (mul_22_8_n_396 ^ mul_22_8_n_387)));
 assign mul_22_8_n_1231 = (mul_22_8_n_653 ^ (mul_22_8_n_396 ^ mul_22_8_n_387));
 assign mul_22_8_n_1223 = ((mul_22_8_n_527 & mul_22_8_n_591) | (mul_22_8_n_518 & (mul_22_8_n_527 ^ mul_22_8_n_591)));
 assign mul_22_8_n_1230 = (mul_22_8_n_518 ^ (mul_22_8_n_527 ^ mul_22_8_n_591));
 assign mul_22_8_n_1220 = ((mul_22_8_n_553 & mul_22_8_n_556) | (mul_22_8_n_699 & (mul_22_8_n_553 ^ mul_22_8_n_556)));
 assign mul_22_8_n_1229 = (mul_22_8_n_699 ^ (mul_22_8_n_553 ^ mul_22_8_n_556));
 assign mul_22_8_n_1218 = ((mul_22_8_n_1232 & mul_22_8_n_1233) | (mul_22_8_n_1231 & (mul_22_8_n_1232
    ^ mul_22_8_n_1233)));
 assign mul_22_8_n_1227 = (mul_22_8_n_1231 ^ (mul_22_8_n_1232 ^ mul_22_8_n_1233));
 assign mul_22_8_n_1216 = ((mul_22_8_n_1229 & mul_22_8_n_1230) | (mul_22_8_n_1228 & (mul_22_8_n_1229
    ^ mul_22_8_n_1230)));
 assign mul_22_8_n_1226 = (mul_22_8_n_1228 ^ (mul_22_8_n_1229 ^ mul_22_8_n_1230));
 assign mul_22_8_n_1300 = ((mul_22_8_n_1226 & mul_22_8_n_1227) | (mul_22_8_n_1225 & (mul_22_8_n_1226
    ^ mul_22_8_n_1227)));
 assign mul_22_8_n_1275 = (mul_22_8_n_1225 ^ (mul_22_8_n_1226 ^ mul_22_8_n_1227));
 assign mul_22_8_n_1214 = ((mul_22_8_n_626 & mul_22_8_n_540) | (mul_22_8_n_536 & (mul_22_8_n_626 ^ mul_22_8_n_540)));
 assign mul_22_8_n_1221 = (mul_22_8_n_536 ^ (mul_22_8_n_626 ^ mul_22_8_n_540));
 assign mul_22_8_n_1213 = ((mul_22_8_n_516 & mul_22_8_n_531) | (mul_22_8_n_528 & (mul_22_8_n_516 ^ mul_22_8_n_531)));
 assign mul_22_8_n_1222 = (mul_22_8_n_528 ^ (mul_22_8_n_516 ^ mul_22_8_n_531));
 assign mul_22_8_n_1209 = ((mul_22_8_n_701 & mul_22_8_n_523) | (mul_22_8_n_1224 & (mul_22_8_n_701 ^ mul_22_8_n_523)));
 assign mul_22_8_n_1219 = (mul_22_8_n_1224 ^ (mul_22_8_n_701 ^ mul_22_8_n_523));
 assign mul_22_8_n_1207 = ((mul_22_8_n_1222 & mul_22_8_n_1223) | (mul_22_8_n_1221 & (mul_22_8_n_1222
    ^ mul_22_8_n_1223)));
 assign mul_22_8_n_1217 = (mul_22_8_n_1221 ^ (mul_22_8_n_1222 ^ mul_22_8_n_1223));
 assign mul_22_8_n_1205 = ((mul_22_8_n_1219 & mul_22_8_n_1220) | (mul_22_8_n_1218 & (mul_22_8_n_1219
    ^ mul_22_8_n_1220)));
 assign mul_22_8_n_1215 = (mul_22_8_n_1218 ^ (mul_22_8_n_1219 ^ mul_22_8_n_1220));
 assign mul_22_8_n_1301 = ((mul_22_8_n_1216 & mul_22_8_n_1217) | (mul_22_8_n_1215 & (mul_22_8_n_1216
    ^ mul_22_8_n_1217)));
 assign mul_22_8_n_1276 = (mul_22_8_n_1215 ^ (mul_22_8_n_1216 ^ mul_22_8_n_1217));
 assign mul_22_8_n_1203 = ((mul_22_8_n_403 & mul_22_8_n_381) | (mul_22_8_n_580 & (mul_22_8_n_403 ^ mul_22_8_n_381)));
 assign mul_22_8_n_1211 = (mul_22_8_n_580 ^ (mul_22_8_n_403 ^ mul_22_8_n_381));
 assign mul_22_8_n_1201 = ((mul_22_8_n_503 & mul_22_8_n_446) | (mul_22_8_n_501 & (mul_22_8_n_503 ^ mul_22_8_n_446)));
 assign mul_22_8_n_1210 = (mul_22_8_n_501 ^ (mul_22_8_n_503 ^ mul_22_8_n_446));
 assign mul_22_8_n_1202 = ((mul_22_8_n_496 & mul_22_8_n_515) | (mul_22_8_n_495 & (mul_22_8_n_496 ^ mul_22_8_n_515)));
 assign mul_22_8_n_1212 = (mul_22_8_n_495 ^ (mul_22_8_n_496 ^ mul_22_8_n_515));
 assign mul_22_8_n_1197 = ((mul_22_8_n_1214 & mul_22_8_n_696) | (mul_22_8_n_1213 & (mul_22_8_n_1214 ^
    mul_22_8_n_696)));
 assign mul_22_8_n_1208 = (mul_22_8_n_1213 ^ (mul_22_8_n_1214 ^ mul_22_8_n_696));
 assign mul_22_8_n_1195 = ((mul_22_8_n_1211 & mul_22_8_n_1212) | (mul_22_8_n_1210 & (mul_22_8_n_1211
    ^ mul_22_8_n_1212)));
 assign mul_22_8_n_1206 = (mul_22_8_n_1210 ^ (mul_22_8_n_1211 ^ mul_22_8_n_1212));
 assign mul_22_8_n_1193 = ((mul_22_8_n_1208 & mul_22_8_n_1209) | (mul_22_8_n_1207 & (mul_22_8_n_1208
    ^ mul_22_8_n_1209)));
 assign mul_22_8_n_1204 = (mul_22_8_n_1207 ^ (mul_22_8_n_1208 ^ mul_22_8_n_1209));
 assign mul_22_8_n_1302 = ((mul_22_8_n_1205 & mul_22_8_n_1206) | (mul_22_8_n_1204 & (mul_22_8_n_1205
    ^ mul_22_8_n_1206)));
 assign mul_22_8_n_1277 = (mul_22_8_n_1204 ^ (mul_22_8_n_1205 ^ mul_22_8_n_1206));
 assign mul_22_8_n_1191 = ((mul_22_8_n_481 & mul_22_8_n_483) | (mul_22_8_n_627 & (mul_22_8_n_481 ^ mul_22_8_n_483)));
 assign mul_22_8_n_1200 = (mul_22_8_n_627 ^ (mul_22_8_n_481 ^ mul_22_8_n_483));
 assign mul_22_8_n_1190 = ((mul_22_8_n_474 & mul_22_8_n_476) | (mul_22_8_n_453 & (mul_22_8_n_474 ^ mul_22_8_n_476)));
 assign mul_22_8_n_1199 = (mul_22_8_n_453 ^ (mul_22_8_n_474 ^ mul_22_8_n_476));
 assign mul_22_8_n_1186 = ((mul_22_8_n_470 & mul_22_8_n_472) | (mul_22_8_n_700 & (mul_22_8_n_470 ^ mul_22_8_n_472)));
 assign mul_22_8_n_1198 = (mul_22_8_n_700 ^ (mul_22_8_n_470 ^ mul_22_8_n_472));
 assign mul_22_8_n_1184 = ((mul_22_8_n_1202 & mul_22_8_n_1203) | (mul_22_8_n_1201 & (mul_22_8_n_1202
    ^ mul_22_8_n_1203)));
 assign mul_22_8_n_1196 = (mul_22_8_n_1201 ^ (mul_22_8_n_1202 ^ mul_22_8_n_1203));
 assign mul_22_8_n_1183 = ((mul_22_8_n_1199 & mul_22_8_n_1200) | (mul_22_8_n_1198 & (mul_22_8_n_1199
    ^ mul_22_8_n_1200)));
 assign mul_22_8_n_1194 = (mul_22_8_n_1198 ^ (mul_22_8_n_1199 ^ mul_22_8_n_1200));
 assign mul_22_8_n_1180 = ((mul_22_8_n_1196 & mul_22_8_n_1197) | (mul_22_8_n_1195 & (mul_22_8_n_1196
    ^ mul_22_8_n_1197)));
 assign mul_22_8_n_1192 = (mul_22_8_n_1195 ^ (mul_22_8_n_1196 ^ mul_22_8_n_1197));
 assign mul_22_8_n_1303 = ((mul_22_8_n_1193 & mul_22_8_n_1194) | (mul_22_8_n_1192 & (mul_22_8_n_1193
    ^ mul_22_8_n_1194)));
 assign mul_22_8_n_1278 = (mul_22_8_n_1192 ^ (mul_22_8_n_1193 ^ mul_22_8_n_1194));
 assign mul_22_8_n_1178 = ((mul_22_8_n_437 & mul_22_8_n_390) | (mul_22_8_n_593 & (mul_22_8_n_437 ^ mul_22_8_n_390)));
 assign mul_22_8_n_1188 = (mul_22_8_n_593 ^ (mul_22_8_n_437 ^ mul_22_8_n_390));
 assign mul_22_8_n_1177 = ((mul_22_8_n_451 & mul_22_8_n_662) | (mul_22_8_n_450 & (mul_22_8_n_451 ^ mul_22_8_n_662)));
 assign mul_22_8_n_1187 = (mul_22_8_n_450 ^ (mul_22_8_n_451 ^ mul_22_8_n_662));
 assign mul_22_8_n_1176 = ((mul_22_8_n_445 & mul_22_8_n_459) | (mul_22_8_n_441 & (mul_22_8_n_445 ^ mul_22_8_n_459)));
 assign mul_22_8_n_1189 = (mul_22_8_n_441 ^ (mul_22_8_n_445 ^ mul_22_8_n_459));
 assign mul_22_8_n_1172 = ((mul_22_8_n_697 & mul_22_8_n_572) | (mul_22_8_n_1191 & (mul_22_8_n_697 ^ mul_22_8_n_572)));
 assign mul_22_8_n_1185 = (mul_22_8_n_1191 ^ (mul_22_8_n_697 ^ mul_22_8_n_572));
 assign mul_22_8_n_1170 = ((mul_22_8_n_1189 & mul_22_8_n_1190) | (mul_22_8_n_1188 & (mul_22_8_n_1189
    ^ mul_22_8_n_1190)));
 assign mul_22_8_n_1182 = (mul_22_8_n_1188 ^ (mul_22_8_n_1189 ^ mul_22_8_n_1190));
 assign mul_22_8_n_1168 = ((mul_22_8_n_1186 & mul_22_8_n_1187) | (mul_22_8_n_1185 & (mul_22_8_n_1186
    ^ mul_22_8_n_1187)));
 assign mul_22_8_n_1181 = (mul_22_8_n_1185 ^ (mul_22_8_n_1186 ^ mul_22_8_n_1187));
 assign mul_22_8_n_1166 = ((mul_22_8_n_1183 & mul_22_8_n_1184) | (mul_22_8_n_1182 & (mul_22_8_n_1183
    ^ mul_22_8_n_1184)));
 assign mul_22_8_n_1179 = (mul_22_8_n_1182 ^ (mul_22_8_n_1183 ^ mul_22_8_n_1184));
 assign mul_22_8_n_1304 = ((mul_22_8_n_1180 & mul_22_8_n_1181) | (mul_22_8_n_1179 & (mul_22_8_n_1180
    ^ mul_22_8_n_1181)));
 assign mul_22_8_n_1279 = (mul_22_8_n_1179 ^ (mul_22_8_n_1180 ^ mul_22_8_n_1181));
 assign mul_22_8_n_1164 = ((mul_22_8_n_614 & mul_22_8_n_471) | (mul_22_8_n_612 & (mul_22_8_n_614 ^ mul_22_8_n_471)));
 assign mul_22_8_n_1174 = (mul_22_8_n_612 ^ (mul_22_8_n_614 ^ mul_22_8_n_471));
 assign mul_22_8_n_1162 = ((mul_22_8_n_628 & mul_22_8_n_609) | (mul_22_8_n_584 & (mul_22_8_n_628 ^ mul_22_8_n_609)));
 assign mul_22_8_n_1173 = (mul_22_8_n_584 ^ (mul_22_8_n_628 ^ mul_22_8_n_609));
 assign mul_22_8_n_1163 = ((mul_22_8_n_657 & mul_22_8_n_600) | (mul_22_8_n_596 & (mul_22_8_n_657 ^ mul_22_8_n_600)));
 assign mul_22_8_n_1175 = (mul_22_8_n_596 ^ (mul_22_8_n_657 ^ mul_22_8_n_600));
 assign mul_22_8_n_1157 = ((mul_22_8_n_1178 & mul_22_8_n_702) | (mul_22_8_n_1177 & (mul_22_8_n_1178 ^
    mul_22_8_n_702)));
 assign mul_22_8_n_1171 = (mul_22_8_n_1177 ^ (mul_22_8_n_1178 ^ mul_22_8_n_702));
 assign mul_22_8_n_1156 = ((mul_22_8_n_1175 & mul_22_8_n_1176) | (mul_22_8_n_1174 & (mul_22_8_n_1175
    ^ mul_22_8_n_1176)));
 assign mul_22_8_n_1169 = (mul_22_8_n_1174 ^ (mul_22_8_n_1175 ^ mul_22_8_n_1176));
 assign mul_22_8_n_1152 = ((mul_22_8_n_1172 & mul_22_8_n_1173) | (mul_22_8_n_1171 & (mul_22_8_n_1172
    ^ mul_22_8_n_1173)));
 assign mul_22_8_n_1167 = (mul_22_8_n_1171 ^ (mul_22_8_n_1172 ^ mul_22_8_n_1173));
 assign mul_22_8_n_1151 = ((mul_22_8_n_1169 & mul_22_8_n_1170) | (mul_22_8_n_1168 & (mul_22_8_n_1169
    ^ mul_22_8_n_1170)));
 assign mul_22_8_n_1165 = (mul_22_8_n_1168 ^ (mul_22_8_n_1169 ^ mul_22_8_n_1170));
 assign mul_22_8_n_1305 = ((mul_22_8_n_1166 & mul_22_8_n_1167) | (mul_22_8_n_1165 & (mul_22_8_n_1166
    ^ mul_22_8_n_1167)));
 assign mul_22_8_n_1280 = (mul_22_8_n_1165 ^ (mul_22_8_n_1166 ^ mul_22_8_n_1167));
 assign mul_22_8_n_1148 = ((mul_22_8_n_409 & mul_22_8_n_389) | (mul_22_8_n_466 & (mul_22_8_n_409 ^ mul_22_8_n_389)));
 assign mul_22_8_n_1161 = (mul_22_8_n_466 ^ (mul_22_8_n_409 ^ mul_22_8_n_389));
 assign mul_22_8_n_1149 = ((mul_22_8_n_574 & mul_22_8_n_520) | (mul_22_8_n_573 & (mul_22_8_n_574 ^ mul_22_8_n_520)));
 assign mul_22_8_n_1160 = (mul_22_8_n_573 ^ (mul_22_8_n_574 ^ mul_22_8_n_520));
 assign mul_22_8_n_1147 = ((mul_22_8_n_604 & mul_22_8_n_585) | (mul_22_8_n_449 & (mul_22_8_n_604 ^ mul_22_8_n_585)));
 assign mul_22_8_n_1159 = (mul_22_8_n_449 ^ (mul_22_8_n_604 ^ mul_22_8_n_585));
 assign mul_22_8_n_1143 = ((mul_22_8_n_454 & mul_22_8_n_569) | (mul_22_8_n_698 & (mul_22_8_n_454 ^ mul_22_8_n_569)));
 assign mul_22_8_n_1158 = (mul_22_8_n_698 ^ (mul_22_8_n_454 ^ mul_22_8_n_569));
 assign mul_22_8_n_1142 = ((mul_22_8_n_1163 & mul_22_8_n_1164) | (mul_22_8_n_1162 & (mul_22_8_n_1163
    ^ mul_22_8_n_1164)));
 assign mul_22_8_n_1155 = (mul_22_8_n_1162 ^ (mul_22_8_n_1163 ^ mul_22_8_n_1164));
 assign mul_22_8_n_1139 = ((mul_22_8_n_1160 & mul_22_8_n_1161) | (mul_22_8_n_1159 & (mul_22_8_n_1160
    ^ mul_22_8_n_1161)));
 assign mul_22_8_n_1154 = (mul_22_8_n_1159 ^ (mul_22_8_n_1160 ^ mul_22_8_n_1161));
 assign mul_22_8_n_1136 = ((mul_22_8_n_1157 & mul_22_8_n_1158) | (mul_22_8_n_1156 & (mul_22_8_n_1157
    ^ mul_22_8_n_1158)));
 assign mul_22_8_n_1153 = (mul_22_8_n_1156 ^ (mul_22_8_n_1157 ^ mul_22_8_n_1158));
 assign mul_22_8_n_1134 = ((mul_22_8_n_1154 & mul_22_8_n_1155) | (mul_22_8_n_1153 & (mul_22_8_n_1154
    ^ mul_22_8_n_1155)));
 assign mul_22_8_n_1150 = (mul_22_8_n_1153 ^ (mul_22_8_n_1154 ^ mul_22_8_n_1155));
 assign mul_22_8_n_1306 = ((mul_22_8_n_1151 & mul_22_8_n_1152) | (mul_22_8_n_1150 & (mul_22_8_n_1151
    ^ mul_22_8_n_1152)));
 assign mul_22_8_n_1281 = (mul_22_8_n_1150 ^ (mul_22_8_n_1151 ^ mul_22_8_n_1152));
 assign mul_22_8_n_1131 = ((mul_22_8_n_533 & mul_22_8_n_469) | (mul_22_8_n_491 & (mul_22_8_n_533 ^ mul_22_8_n_469)));
 assign mul_22_8_n_1145 = (mul_22_8_n_491 ^ (mul_22_8_n_533 ^ mul_22_8_n_469));
 assign mul_22_8_n_1132 = ((mul_22_8_n_509 & mul_22_8_n_664) | (mul_22_8_n_630 & (mul_22_8_n_509 ^ mul_22_8_n_664)));
 assign mul_22_8_n_1144 = (mul_22_8_n_630 ^ (mul_22_8_n_509 ^ mul_22_8_n_664));
 assign mul_22_8_n_1133 = ((mul_22_8_n_468 & mul_22_8_n_404) | (mul_22_8_n_568 & (mul_22_8_n_468 ^ mul_22_8_n_404)));
 assign mul_22_8_n_1146 = (mul_22_8_n_568 ^ (mul_22_8_n_468 ^ mul_22_8_n_404));
 assign mul_22_8_n_1126 = ((mul_22_8_n_713 & mul_22_8_n_660) | (mul_22_8_n_1149 & (mul_22_8_n_713 ^ mul_22_8_n_660)));
 assign mul_22_8_n_1141 = (mul_22_8_n_1149 ^ (mul_22_8_n_713 ^ mul_22_8_n_660));
 assign mul_22_8_n_1125 = ((mul_22_8_n_1147 & mul_22_8_n_1148) | (mul_22_8_n_1146 & (mul_22_8_n_1147
    ^ mul_22_8_n_1148)));
 assign mul_22_8_n_1140 = (mul_22_8_n_1146 ^ (mul_22_8_n_1147 ^ mul_22_8_n_1148));
 assign mul_22_8_n_1123 = ((mul_22_8_n_1144 & mul_22_8_n_1145) | (mul_22_8_n_1143 & (mul_22_8_n_1144
    ^ mul_22_8_n_1145)));
 assign mul_22_8_n_1138 = (mul_22_8_n_1143 ^ (mul_22_8_n_1144 ^ mul_22_8_n_1145));
 assign mul_22_8_n_1120 = ((mul_22_8_n_1141 & mul_22_8_n_1142) | (mul_22_8_n_1140 & (mul_22_8_n_1141
    ^ mul_22_8_n_1142)));
 assign mul_22_8_n_1137 = (mul_22_8_n_1140 ^ (mul_22_8_n_1141 ^ mul_22_8_n_1142));
 assign mul_22_8_n_1117 = ((mul_22_8_n_1138 & mul_22_8_n_1139) | (mul_22_8_n_1137 & (mul_22_8_n_1138
    ^ mul_22_8_n_1139)));
 assign mul_22_8_n_1135 = (mul_22_8_n_1137 ^ (mul_22_8_n_1138 ^ mul_22_8_n_1139));
 assign mul_22_8_n_1307 = ((n_57 & n_35) | (n_77 & (n_57 ^ n_35)));
 assign mul_22_8_n_1282 = (n_77 ^ (n_57 ^ n_35));
 assign mul_22_8_n_1114 = ((mul_22_8_n_555 & mul_22_8_n_383) | (mul_22_8_n_554 & (mul_22_8_n_555 ^ mul_22_8_n_383)));
 assign mul_22_8_n_1127 = (mul_22_8_n_554 ^ (mul_22_8_n_555 ^ mul_22_8_n_383));
 assign mul_22_8_n_1113 = ((mul_22_8_n_550 & mul_22_8_n_552) | (mul_22_8_n_549 & (mul_22_8_n_550 ^ mul_22_8_n_552)));
 assign mul_22_8_n_1129 = (mul_22_8_n_549 ^ (mul_22_8_n_550 ^ mul_22_8_n_552));
 assign mul_22_8_n_1116 = ((mul_22_8_n_547 & mul_22_8_n_548) | (mul_22_8_n_398 & (mul_22_8_n_547 ^ mul_22_8_n_548)));
 assign mul_22_8_n_1128 = (mul_22_8_n_398 ^ (mul_22_8_n_547 ^ mul_22_8_n_548));
 assign mul_22_8_n_1115 = ((mul_22_8_n_544 & mul_22_8_n_545) | (mul_22_8_n_543 & (mul_22_8_n_544 ^ mul_22_8_n_545)));
 assign mul_22_8_n_1130 = (mul_22_8_n_543 ^ (mul_22_8_n_544 ^ mul_22_8_n_545));
 assign mul_22_8_n_1108 = ((mul_22_8_n_1133 & mul_22_8_n_690) | (mul_22_8_n_1132 & (mul_22_8_n_1133 ^
    mul_22_8_n_690)));
 assign mul_22_8_n_1124 = (mul_22_8_n_1132 ^ (mul_22_8_n_1133 ^ mul_22_8_n_690));
 assign mul_22_8_n_1106 = ((mul_22_8_n_1130 & mul_22_8_n_1131) | (mul_22_8_n_1129 & (mul_22_8_n_1130
    ^ mul_22_8_n_1131)));
 assign mul_22_8_n_1122 = (mul_22_8_n_1129 ^ (mul_22_8_n_1130 ^ mul_22_8_n_1131));
 assign mul_22_8_n_1103 = ((mul_22_8_n_1127 & mul_22_8_n_1128) | (mul_22_8_n_1126 & (mul_22_8_n_1127
    ^ mul_22_8_n_1128)));
 assign mul_22_8_n_1121 = (mul_22_8_n_1126 ^ (mul_22_8_n_1127 ^ mul_22_8_n_1128));
 assign mul_22_8_n_1101 = ((mul_22_8_n_1124 & mul_22_8_n_1125) | (mul_22_8_n_1123 & (mul_22_8_n_1124
    ^ mul_22_8_n_1125)));
 assign mul_22_8_n_1119 = (mul_22_8_n_1123 ^ (mul_22_8_n_1124 ^ mul_22_8_n_1125));
 assign mul_22_8_n_1100 = ((mul_22_8_n_1121 & mul_22_8_n_1122) | (mul_22_8_n_1120 & (mul_22_8_n_1121
    ^ mul_22_8_n_1122)));
 assign mul_22_8_n_1118 = (mul_22_8_n_1120 ^ (mul_22_8_n_1121 ^ mul_22_8_n_1122));
 assign mul_22_8_n_1308 = ((mul_22_8_n_1118 & mul_22_8_n_1119) | (mul_22_8_n_1117 & (mul_22_8_n_1118
    ^ mul_22_8_n_1119)));
 assign mul_22_8_n_1283 = (mul_22_8_n_1117 ^ (mul_22_8_n_1118 ^ mul_22_8_n_1119));
 assign mul_22_8_n_1096 = ((mul_22_8_n_530 & mul_22_8_n_532) | (mul_22_8_n_529 & (mul_22_8_n_530 ^ mul_22_8_n_532)));
 assign mul_22_8_n_1110 = (mul_22_8_n_529 ^ (mul_22_8_n_530 ^ mul_22_8_n_532));
 assign mul_22_8_n_1098 = ((mul_22_8_n_525 & mul_22_8_n_546) | (mul_22_8_n_524 & (mul_22_8_n_525 ^ mul_22_8_n_546)));
 assign mul_22_8_n_1111 = (mul_22_8_n_524 ^ (mul_22_8_n_525 ^ mul_22_8_n_546));
 assign mul_22_8_n_1097 = ((mul_22_8_n_522 & mul_22_8_n_395) | (mul_22_8_n_632 & (mul_22_8_n_522 ^ mul_22_8_n_395)));
 assign mul_22_8_n_1112 = (mul_22_8_n_632 ^ (mul_22_8_n_522 ^ mul_22_8_n_395));
 assign mul_22_8_n_1091 = ((mul_22_8_n_500 & mul_22_8_n_521) | (mul_22_8_n_712 & (mul_22_8_n_500 ^ mul_22_8_n_521)));
 assign mul_22_8_n_1109 = (mul_22_8_n_712 ^ (mul_22_8_n_500 ^ mul_22_8_n_521));
 assign mul_22_8_n_1090 = ((mul_22_8_n_1115 & mul_22_8_n_1116) | (mul_22_8_n_1114 & (mul_22_8_n_1115
    ^ mul_22_8_n_1116)));
 assign mul_22_8_n_1107 = (mul_22_8_n_1114 ^ (mul_22_8_n_1115 ^ mul_22_8_n_1116));
 assign mul_22_8_n_1087 = ((mul_22_8_n_1112 & mul_22_8_n_1113) | (mul_22_8_n_1111 & (mul_22_8_n_1112
    ^ mul_22_8_n_1113)));
 assign mul_22_8_n_1105 = (mul_22_8_n_1111 ^ (mul_22_8_n_1112 ^ mul_22_8_n_1113));
 assign mul_22_8_n_1085 = ((mul_22_8_n_1109 & mul_22_8_n_1110) | (mul_22_8_n_1108 & (mul_22_8_n_1109
    ^ mul_22_8_n_1110)));
 assign mul_22_8_n_1104 = (mul_22_8_n_1108 ^ (mul_22_8_n_1109 ^ mul_22_8_n_1110));
 assign mul_22_8_n_1083 = ((mul_22_8_n_1106 & mul_22_8_n_1107) | (mul_22_8_n_1105 & (mul_22_8_n_1106
    ^ mul_22_8_n_1107)));
 assign mul_22_8_n_1102 = (mul_22_8_n_1105 ^ (mul_22_8_n_1106 ^ mul_22_8_n_1107));
 assign mul_22_8_n_1080 = ((mul_22_8_n_1103 & mul_22_8_n_1104) | (mul_22_8_n_1102 & (mul_22_8_n_1103
    ^ mul_22_8_n_1104)));
 assign mul_22_8_n_1099 = (mul_22_8_n_1102 ^ (mul_22_8_n_1103 ^ mul_22_8_n_1104));
 assign mul_22_8_n_1309 = ((n_74 & n_58) | (n_80 & (n_74 ^ n_58)));
 assign mul_22_8_n_1284 = (n_80 ^ (n_74 ^ n_58));
 assign mul_22_8_n_1076 = ((mul_22_8_n_508 & mul_22_8_n_393) | (mul_22_8_n_507 & (mul_22_8_n_508 ^ mul_22_8_n_393)));
 assign mul_22_8_n_1093 = (mul_22_8_n_507 ^ (mul_22_8_n_508 ^ mul_22_8_n_393));
 assign mul_22_8_n_1079 = ((mul_22_8_n_594 & mul_22_8_n_588) | (mul_22_8_n_603 & (mul_22_8_n_594 ^ mul_22_8_n_588)));
 assign mul_22_8_n_1092 = (mul_22_8_n_603 ^ (mul_22_8_n_594 ^ mul_22_8_n_588));
 assign mul_22_8_n_1078 = ((mul_22_8_n_502 & mul_22_8_n_504) | (mul_22_8_n_408 & (mul_22_8_n_502 ^ mul_22_8_n_504)));
 assign mul_22_8_n_1094 = (mul_22_8_n_408 ^ (mul_22_8_n_502 ^ mul_22_8_n_504));
 assign mul_22_8_n_1077 = ((mul_22_8_n_498 & mul_22_8_n_499) | (mul_22_8_n_537 & (mul_22_8_n_498 ^ mul_22_8_n_499)));
 assign mul_22_8_n_1095 = (mul_22_8_n_537 ^ (mul_22_8_n_498 ^ mul_22_8_n_499));
 assign mul_22_8_n_1071 = ((mul_22_8_n_688 & mul_22_8_n_497) | (mul_22_8_n_1098 & (mul_22_8_n_688 ^ mul_22_8_n_497)));
 assign mul_22_8_n_1089 = (mul_22_8_n_1098 ^ (mul_22_8_n_688 ^ mul_22_8_n_497));
 assign mul_22_8_n_1068 = ((mul_22_8_n_1096 & mul_22_8_n_1097) | (mul_22_8_n_1095 & (mul_22_8_n_1096
    ^ mul_22_8_n_1097)));
 assign mul_22_8_n_1088 = (mul_22_8_n_1095 ^ (mul_22_8_n_1096 ^ mul_22_8_n_1097));
 assign mul_22_8_n_1069 = ((mul_22_8_n_1093 & mul_22_8_n_1094) | (mul_22_8_n_1092 & (mul_22_8_n_1093
    ^ mul_22_8_n_1094)));
 assign mul_22_8_n_1086 = (mul_22_8_n_1092 ^ (mul_22_8_n_1093 ^ mul_22_8_n_1094));
 assign mul_22_8_n_1065 = ((mul_22_8_n_1090 & mul_22_8_n_1091) | (mul_22_8_n_1089 & (mul_22_8_n_1090
    ^ mul_22_8_n_1091)));
 assign mul_22_8_n_1084 = (mul_22_8_n_1089 ^ (mul_22_8_n_1090 ^ mul_22_8_n_1091));
 assign mul_22_8_n_1064 = ((mul_22_8_n_1087 & mul_22_8_n_1088) | (mul_22_8_n_1086 & (mul_22_8_n_1087
    ^ mul_22_8_n_1088)));
 assign mul_22_8_n_1082 = (mul_22_8_n_1086 ^ (mul_22_8_n_1087 ^ mul_22_8_n_1088));
 assign mul_22_8_n_1061 = ((mul_22_8_n_1084 & mul_22_8_n_1085) | (mul_22_8_n_1083 & (mul_22_8_n_1084
    ^ mul_22_8_n_1085)));
 assign mul_22_8_n_1081 = (mul_22_8_n_1083 ^ (mul_22_8_n_1084 ^ mul_22_8_n_1085));
 assign mul_22_8_n_1310 = ((mul_22_8_n_1081 & mul_22_8_n_1082) | (mul_22_8_n_1080 & (mul_22_8_n_1081
    ^ mul_22_8_n_1082)));
 assign mul_22_8_n_1285 = (mul_22_8_n_1080 ^ (mul_22_8_n_1081 ^ mul_22_8_n_1082));
 assign mul_22_8_n_1059 = ((mul_22_8_n_487 & mul_22_8_n_488) | (mul_22_8_n_473 & (mul_22_8_n_487 ^ mul_22_8_n_488)));
 assign mul_22_8_n_1074 = (mul_22_8_n_473 ^ (mul_22_8_n_487 ^ mul_22_8_n_488));
 assign mul_22_8_n_1058 = ((mul_22_8_n_484 & mul_22_8_n_485) | (mul_22_8_n_514 & (mul_22_8_n_484 ^ mul_22_8_n_485)));
 assign mul_22_8_n_1073 = (mul_22_8_n_514 ^ (mul_22_8_n_484 ^ mul_22_8_n_485));
 assign mul_22_8_n_1057 = ((mul_22_8_n_482 & mul_22_8_n_406) | (mul_22_8_n_480 & (mul_22_8_n_482 ^ mul_22_8_n_406)));
 assign mul_22_8_n_1072 = (mul_22_8_n_480 ^ (mul_22_8_n_482 ^ mul_22_8_n_406));
 assign mul_22_8_n_1056 = ((mul_22_8_n_479 & mul_22_8_n_634) | (mul_22_8_n_478 & (mul_22_8_n_479 ^ mul_22_8_n_634)));
 assign mul_22_8_n_1075 = (mul_22_8_n_478 ^ (mul_22_8_n_479 ^ mul_22_8_n_634));
 assign mul_22_8_n_1050 = ((mul_22_8_n_1079 & mul_22_8_n_708) | (mul_22_8_n_1078 & (mul_22_8_n_1079 ^
    mul_22_8_n_708)));
 assign mul_22_8_n_1067 = (mul_22_8_n_1078 ^ (mul_22_8_n_1079 ^ mul_22_8_n_708));
 assign mul_22_8_n_1049 = ((mul_22_8_n_1076 & mul_22_8_n_1077) | (mul_22_8_n_1075 & (mul_22_8_n_1076
    ^ mul_22_8_n_1077)));
 assign mul_22_8_n_1070 = (mul_22_8_n_1075 ^ (mul_22_8_n_1076 ^ mul_22_8_n_1077));
 assign mul_22_8_n_1048 = ((mul_22_8_n_1073 & mul_22_8_n_1074) | (mul_22_8_n_1072 & (mul_22_8_n_1073
    ^ mul_22_8_n_1074)));
 assign mul_22_8_n_1066 = (mul_22_8_n_1072 ^ (mul_22_8_n_1073 ^ mul_22_8_n_1074));
 assign mul_22_8_n_1044 = ((mul_22_8_n_1070 & mul_22_8_n_1071) | (mul_22_8_n_1069 & (mul_22_8_n_1070
    ^ mul_22_8_n_1071)));
 assign mul_22_8_n_1063 = (mul_22_8_n_1069 ^ (mul_22_8_n_1070 ^ mul_22_8_n_1071));
 assign mul_22_8_n_1042 = ((mul_22_8_n_1067 & mul_22_8_n_1068) | (mul_22_8_n_1066 & (mul_22_8_n_1067
    ^ mul_22_8_n_1068)));
 assign mul_22_8_n_1062 = (mul_22_8_n_1066 ^ (mul_22_8_n_1067 ^ mul_22_8_n_1068));
 assign mul_22_8_n_1040 = ((mul_22_8_n_1064 & mul_22_8_n_1065) | (mul_22_8_n_1063 & (mul_22_8_n_1064
    ^ mul_22_8_n_1065)));
 assign mul_22_8_n_1060 = (mul_22_8_n_1063 ^ (mul_22_8_n_1064 ^ mul_22_8_n_1065));
 assign mul_22_8_n_1311 = ((n_40 & n_70) | (n_59 & (n_40 ^ n_70)));
 assign mul_22_8_n_1286 = (n_59 ^ (n_40 ^ n_70));
 assign mul_22_8_n_1038 = ((mul_22_8_n_467 & mul_22_8_n_380) | (mul_22_8_n_475 & (mul_22_8_n_467 ^ mul_22_8_n_380)));
 assign mul_22_8_n_1055 = (mul_22_8_n_475 ^ (mul_22_8_n_467 ^ mul_22_8_n_380));
 assign mul_22_8_n_1037 = ((mul_22_8_n_464 & mul_22_8_n_517) | (mul_22_8_n_463 & (mul_22_8_n_464 ^ mul_22_8_n_517)));
 assign mul_22_8_n_1053 = (mul_22_8_n_463 ^ (mul_22_8_n_464 ^ mul_22_8_n_517));
 assign mul_22_8_n_1036 = ((mul_22_8_n_460 & mul_22_8_n_461) | (mul_22_8_n_407 & (mul_22_8_n_460 ^ mul_22_8_n_461)));
 assign mul_22_8_n_1054 = (mul_22_8_n_407 ^ (mul_22_8_n_460 ^ mul_22_8_n_461));
 assign mul_22_8_n_1035 = ((mul_22_8_n_456 & mul_22_8_n_457) | (mul_22_8_n_661 & (mul_22_8_n_456 ^ mul_22_8_n_457)));
 assign mul_22_8_n_1052 = (mul_22_8_n_661 ^ (mul_22_8_n_456 ^ mul_22_8_n_457));
 assign mul_22_8_n_1030 = ((mul_22_8_n_564 & mul_22_8_n_455) | (mul_22_8_n_689 & (mul_22_8_n_564 ^ mul_22_8_n_455)));
 assign mul_22_8_n_1051 = (mul_22_8_n_689 ^ (mul_22_8_n_564 ^ mul_22_8_n_455));
 assign mul_22_8_n_1028 = ((mul_22_8_n_1058 & mul_22_8_n_1059) | (mul_22_8_n_1057 & (mul_22_8_n_1058
    ^ mul_22_8_n_1059)));
 assign mul_22_8_n_1047 = (mul_22_8_n_1057 ^ (mul_22_8_n_1058 ^ mul_22_8_n_1059));
 assign mul_22_8_n_1027 = ((mul_22_8_n_1055 & mul_22_8_n_1056) | (mul_22_8_n_1054 & (mul_22_8_n_1055
    ^ mul_22_8_n_1056)));
 assign mul_22_8_n_1045 = (mul_22_8_n_1054 ^ (mul_22_8_n_1055 ^ mul_22_8_n_1056));
 assign mul_22_8_n_1025 = ((mul_22_8_n_1052 & mul_22_8_n_1053) | (mul_22_8_n_1051 & (mul_22_8_n_1052
    ^ mul_22_8_n_1053)));
 assign mul_22_8_n_1046 = (mul_22_8_n_1051 ^ (mul_22_8_n_1052 ^ mul_22_8_n_1053));
 assign mul_22_8_n_1022 = ((mul_22_8_n_1049 & mul_22_8_n_1050) | (mul_22_8_n_1048 & (mul_22_8_n_1049
    ^ mul_22_8_n_1050)));
 assign mul_22_8_n_1043 = (mul_22_8_n_1048 ^ (mul_22_8_n_1049 ^ mul_22_8_n_1050));
 assign mul_22_8_n_1021 = ((mul_22_8_n_1046 & mul_22_8_n_1047) | (mul_22_8_n_1045 & (mul_22_8_n_1046
    ^ mul_22_8_n_1047)));
 assign mul_22_8_n_1041 = (mul_22_8_n_1045 ^ (mul_22_8_n_1046 ^ mul_22_8_n_1047));
 assign mul_22_8_n_1018 = ((mul_22_8_n_1043 & mul_22_8_n_1044) | (mul_22_8_n_1042 & (mul_22_8_n_1043
    ^ mul_22_8_n_1044)));
 assign mul_22_8_n_1039 = (mul_22_8_n_1042 ^ (mul_22_8_n_1043 ^ mul_22_8_n_1044));
 assign mul_22_8_n_1312 = ((mul_22_8_n_1040 & mul_22_8_n_1041) | (mul_22_8_n_1039 & (mul_22_8_n_1040
    ^ mul_22_8_n_1041)));
 assign mul_22_8_n_1287 = (mul_22_8_n_1039 ^ (mul_22_8_n_1040 ^ mul_22_8_n_1041));
 assign mul_22_8_n_1016 = ((mul_22_8_n_447 & mul_22_8_n_448) | (mul_22_8_n_465 & (mul_22_8_n_447 ^ mul_22_8_n_448)));
 assign mul_22_8_n_1033 = (mul_22_8_n_465 ^ (mul_22_8_n_447 ^ mul_22_8_n_448));
 assign mul_22_8_n_1015 = ((mul_22_8_n_442 & mul_22_8_n_444) | (mul_22_8_n_506 & (mul_22_8_n_442 ^ mul_22_8_n_444)));
 assign mul_22_8_n_1031 = (mul_22_8_n_506 ^ (mul_22_8_n_442 ^ mul_22_8_n_444));
 assign mul_22_8_n_1013 = ((mul_22_8_n_592 & mul_22_8_n_399) | (mul_22_8_n_654 & (mul_22_8_n_592 ^ mul_22_8_n_399)));
 assign mul_22_8_n_1032 = (mul_22_8_n_654 ^ (mul_22_8_n_592 ^ mul_22_8_n_399));
 assign mul_22_8_n_1014 = ((mul_22_8_n_589 & mul_22_8_n_587) | (mul_22_8_n_637 & (mul_22_8_n_589 ^ mul_22_8_n_587)));
 assign mul_22_8_n_1034 = (mul_22_8_n_637 ^ (mul_22_8_n_589 ^ mul_22_8_n_587));
 assign mul_22_8_n_1006 = ((mul_22_8_n_710 & mul_22_8_n_505) | (mul_22_8_n_1038 & (mul_22_8_n_710 ^ mul_22_8_n_505)));
 assign mul_22_8_n_1029 = (mul_22_8_n_1038 ^ (mul_22_8_n_710 ^ mul_22_8_n_505));
 assign mul_22_8_n_1007 = ((mul_22_8_n_1036 & mul_22_8_n_1037) | (mul_22_8_n_1035 & (mul_22_8_n_1036
    ^ mul_22_8_n_1037)));
 assign mul_22_8_n_1026 = (mul_22_8_n_1035 ^ (mul_22_8_n_1036 ^ mul_22_8_n_1037));
 assign mul_22_8_n_1003 = ((mul_22_8_n_1033 & mul_22_8_n_1034) | (mul_22_8_n_1032 & (mul_22_8_n_1033
    ^ mul_22_8_n_1034)));
 assign mul_22_8_n_1024 = (mul_22_8_n_1032 ^ (mul_22_8_n_1033 ^ mul_22_8_n_1034));
 assign mul_22_8_n_1001 = ((mul_22_8_n_1030 & mul_22_8_n_1031) | (mul_22_8_n_1029 & (mul_22_8_n_1030
    ^ mul_22_8_n_1031)));
 assign mul_22_8_n_1023 = (mul_22_8_n_1029 ^ (mul_22_8_n_1030 ^ mul_22_8_n_1031));
 assign mul_22_8_n_1000 = ((mul_22_8_n_1027 & mul_22_8_n_1028) | (mul_22_8_n_1026 & (mul_22_8_n_1027
    ^ mul_22_8_n_1028)));
 assign mul_22_8_n_1020 = (mul_22_8_n_1026 ^ (mul_22_8_n_1027 ^ mul_22_8_n_1028));
 assign mul_22_8_n_997 = ((mul_22_8_n_1024 & mul_22_8_n_1025) | (mul_22_8_n_1023 & (mul_22_8_n_1024 ^
    mul_22_8_n_1025)));
 assign mul_22_8_n_1019 = (mul_22_8_n_1023 ^ (mul_22_8_n_1024 ^ mul_22_8_n_1025));
 assign mul_22_8_n_995 = ((mul_22_8_n_1021 & mul_22_8_n_1022) | (mul_22_8_n_1020 & (mul_22_8_n_1021 ^
    mul_22_8_n_1022)));
 assign mul_22_8_n_1017 = (mul_22_8_n_1020 ^ (mul_22_8_n_1021 ^ mul_22_8_n_1022));
 assign mul_22_8_n_1313 = ((n_69 & n_23) | (n_43 & (n_69 ^ n_23)));
 assign mul_22_8_n_1288 = (n_43 ^ (n_69 ^ n_23));
 assign mul_22_8_n_992 = ((mul_22_8_n_610 & mul_22_8_n_392) | (mul_22_8_n_659 & (mul_22_8_n_610 ^ mul_22_8_n_392)));
 assign mul_22_8_n_1010 = (mul_22_8_n_659 ^ (mul_22_8_n_610 ^ mul_22_8_n_392));
 assign mul_22_8_n_991 = ((mul_22_8_n_608 & mul_22_8_n_586) | (mul_22_8_n_512 & (mul_22_8_n_608 ^ mul_22_8_n_586)));
 assign mul_22_8_n_1012 = (mul_22_8_n_512 ^ (mul_22_8_n_608 ^ mul_22_8_n_586));
 assign mul_22_8_n_993 = ((mul_22_8_n_606 & mul_22_8_n_607) | (mul_22_8_n_419 & (mul_22_8_n_606 ^ mul_22_8_n_607)));
 assign mul_22_8_n_1009 = (mul_22_8_n_419 ^ (mul_22_8_n_606 ^ mul_22_8_n_607));
 assign mul_22_8_n_990 = ((mul_22_8_n_602 & mul_22_8_n_656) | (mul_22_8_n_601 & (mul_22_8_n_602 ^ mul_22_8_n_656)));
 assign mul_22_8_n_1008 = (mul_22_8_n_601 ^ (mul_22_8_n_602 ^ mul_22_8_n_656));
 assign mul_22_8_n_989 = ((mul_22_8_n_597 & mul_22_8_n_598) | (mul_22_8_n_595 & (mul_22_8_n_597 ^ mul_22_8_n_598)));
 assign mul_22_8_n_1011 = (mul_22_8_n_595 ^ (mul_22_8_n_597 ^ mul_22_8_n_598));
 assign mul_22_8_n_983 = ((mul_22_8_n_1016 & mul_22_8_n_693) | (mul_22_8_n_1015 & (mul_22_8_n_1016 ^
    mul_22_8_n_693)));
 assign mul_22_8_n_1005 = (mul_22_8_n_1015 ^ (mul_22_8_n_1016 ^ mul_22_8_n_693));
 assign mul_22_8_n_980 = ((mul_22_8_n_1013 & mul_22_8_n_1014) | (mul_22_8_n_1012 & (mul_22_8_n_1013 ^
    mul_22_8_n_1014)));
 assign mul_22_8_n_1004 = (mul_22_8_n_1012 ^ (mul_22_8_n_1013 ^ mul_22_8_n_1014));
 assign mul_22_8_n_982 = ((mul_22_8_n_1010 & mul_22_8_n_1011) | (mul_22_8_n_1009 & (mul_22_8_n_1010 ^
    mul_22_8_n_1011)));
 assign mul_22_8_n_1002 = (mul_22_8_n_1009 ^ (mul_22_8_n_1010 ^ mul_22_8_n_1011));
 assign mul_22_8_n_977 = ((mul_22_8_n_1007 & mul_22_8_n_1008) | (mul_22_8_n_1006 & (mul_22_8_n_1007 ^
    mul_22_8_n_1008)));
 assign mul_22_8_n_999 = (mul_22_8_n_1006 ^ (mul_22_8_n_1007 ^ mul_22_8_n_1008));
 assign mul_22_8_n_976 = ((mul_22_8_n_1004 & mul_22_8_n_1005) | (mul_22_8_n_1003 & (mul_22_8_n_1004 ^
    mul_22_8_n_1005)));
 assign mul_22_8_n_998 = (mul_22_8_n_1003 ^ (mul_22_8_n_1004 ^ mul_22_8_n_1005));
 assign mul_22_8_n_972 = ((mul_22_8_n_1001 & mul_22_8_n_1002) | (mul_22_8_n_1000 & (mul_22_8_n_1001 ^
    mul_22_8_n_1002)));
 assign mul_22_8_n_996 = (mul_22_8_n_1000 ^ (mul_22_8_n_1001 ^ mul_22_8_n_1002));
 assign mul_22_8_n_971 = ((mul_22_8_n_998 & mul_22_8_n_999) | (mul_22_8_n_997 & (mul_22_8_n_998 ^ mul_22_8_n_999)));
 assign mul_22_8_n_994 = (mul_22_8_n_997 ^ (mul_22_8_n_998 ^ mul_22_8_n_999));
 assign mul_22_8_n_1314 = ((n_44 & n_84) | (n_55 & (n_44 ^ n_84)));
 assign mul_22_8_n_1289 = (n_55 ^ (n_44 ^ n_84));
 assign mul_22_8_n_969 = ((mul_22_8_n_570 & mul_22_8_n_663) | (mul_22_8_n_452 & (mul_22_8_n_570 ^ mul_22_8_n_663)));
 assign mul_22_8_n_988 = (mul_22_8_n_452 ^ (mul_22_8_n_570 ^ mul_22_8_n_663));
 assign mul_22_8_n_968 = ((mul_22_8_n_583 & mul_22_8_n_489) | (mul_22_8_n_535 & (mul_22_8_n_583 ^ mul_22_8_n_489)));
 assign mul_22_8_n_986 = (mul_22_8_n_535 ^ (mul_22_8_n_583 ^ mul_22_8_n_489));
 assign mul_22_8_n_967 = ((mul_22_8_n_579 & mul_22_8_n_647) | (mul_22_8_n_581 & (mul_22_8_n_579 ^ mul_22_8_n_647)));
 assign mul_22_8_n_985 = (mul_22_8_n_581 ^ (mul_22_8_n_579 ^ mul_22_8_n_647));
 assign mul_22_8_n_966 = ((mul_22_8_n_578 & mul_22_8_n_486) | (mul_22_8_n_538 & (mul_22_8_n_578 ^ mul_22_8_n_486)));
 assign mul_22_8_n_987 = (mul_22_8_n_538 ^ (mul_22_8_n_578 ^ mul_22_8_n_486));
 assign mul_22_8_n_960 = ((mul_22_8_n_640 & mul_22_8_n_575) | (mul_22_8_n_705 & (mul_22_8_n_640 ^ mul_22_8_n_575)));
 assign mul_22_8_n_984 = (mul_22_8_n_705 ^ (mul_22_8_n_640 ^ mul_22_8_n_575));
 assign mul_22_8_n_958 = ((mul_22_8_n_992 & mul_22_8_n_993) | (mul_22_8_n_991 & (mul_22_8_n_992 ^ mul_22_8_n_993)));
 assign mul_22_8_n_981 = (mul_22_8_n_991 ^ (mul_22_8_n_992 ^ mul_22_8_n_993));
 assign mul_22_8_n_955 = ((mul_22_8_n_989 & mul_22_8_n_990) | (mul_22_8_n_988 & (mul_22_8_n_989 ^ mul_22_8_n_990)));
 assign mul_22_8_n_979 = (mul_22_8_n_988 ^ (mul_22_8_n_989 ^ mul_22_8_n_990));
 assign mul_22_8_n_957 = ((mul_22_8_n_986 & mul_22_8_n_987) | (mul_22_8_n_985 & (mul_22_8_n_986 ^ mul_22_8_n_987)));
 assign mul_22_8_n_978 = (mul_22_8_n_985 ^ (mul_22_8_n_986 ^ mul_22_8_n_987));
 assign mul_22_8_n_951 = ((mul_22_8_n_983 & mul_22_8_n_984) | (mul_22_8_n_982 & (mul_22_8_n_983 ^ mul_22_8_n_984)));
 assign mul_22_8_n_975 = (mul_22_8_n_982 ^ (mul_22_8_n_983 ^ mul_22_8_n_984));
 assign mul_22_8_n_952 = ((mul_22_8_n_980 & mul_22_8_n_981) | (mul_22_8_n_979 & (mul_22_8_n_980 ^ mul_22_8_n_981)));
 assign mul_22_8_n_974 = (mul_22_8_n_979 ^ (mul_22_8_n_980 ^ mul_22_8_n_981));
 assign mul_22_8_n_948 = ((mul_22_8_n_977 & mul_22_8_n_978) | (mul_22_8_n_976 & (mul_22_8_n_977 ^ mul_22_8_n_978)));
 assign mul_22_8_n_973 = (mul_22_8_n_976 ^ (mul_22_8_n_977 ^ mul_22_8_n_978));
 assign mul_22_8_n_945 = ((mul_22_8_n_974 & mul_22_8_n_975) | (mul_22_8_n_973 & (mul_22_8_n_974 ^ mul_22_8_n_975)));
 assign mul_22_8_n_970 = (mul_22_8_n_973 ^ (mul_22_8_n_974 ^ mul_22_8_n_975));
 assign mul_22_8_n_1315 = ((n_56 & n_85) | (n_53 & (n_56 ^ n_85)));
 assign mul_22_8_n_1290 = (n_53 ^ (n_56 ^ n_85));
 assign mul_22_8_n_944 = ((mul_22_8_n_420 & mul_22_8_n_382) | (mul_22_8_n_655 & (mul_22_8_n_420 ^ mul_22_8_n_382)));
 assign mul_22_8_n_965 = (mul_22_8_n_655 ^ (mul_22_8_n_420 ^ mul_22_8_n_382));
 assign mul_22_8_n_943 = ((mul_22_8_n_565 & mul_22_8_n_615) | (mul_22_8_n_617 & (mul_22_8_n_565 ^ mul_22_8_n_615)));
 assign mul_22_8_n_961 = (mul_22_8_n_617 ^ (mul_22_8_n_565 ^ mul_22_8_n_615));
 assign mul_22_8_n_942 = ((mul_22_8_n_443 & mul_22_8_n_613) | (mul_22_8_n_511 & (mul_22_8_n_443 ^ mul_22_8_n_613)));
 assign mul_22_8_n_962 = (mul_22_8_n_511 ^ (mul_22_8_n_443 ^ mul_22_8_n_613));
 assign mul_22_8_n_941 = ((mul_22_8_n_648 & mul_22_8_n_526) | (mul_22_8_n_577 & (mul_22_8_n_648 ^ mul_22_8_n_526)));
 assign mul_22_8_n_963 = (mul_22_8_n_577 ^ (mul_22_8_n_648 ^ mul_22_8_n_526));
 assign mul_22_8_n_940 = ((mul_22_8_n_650 & mul_22_8_n_649) | (mul_22_8_n_493 & (mul_22_8_n_650 ^ mul_22_8_n_649)));
 assign mul_22_8_n_964 = (mul_22_8_n_493 ^ (mul_22_8_n_650 ^ mul_22_8_n_649));
 assign mul_22_8_n_933 = ((mul_22_8_n_695 & mul_22_8_n_652) | (mul_22_8_n_969 & (mul_22_8_n_695 ^ mul_22_8_n_652)));
 assign mul_22_8_n_959 = (mul_22_8_n_969 ^ (mul_22_8_n_695 ^ mul_22_8_n_652));
 assign mul_22_8_n_934 = ((mul_22_8_n_967 & mul_22_8_n_968) | (mul_22_8_n_966 & (mul_22_8_n_967 ^ mul_22_8_n_968)));
 assign mul_22_8_n_956 = (mul_22_8_n_966 ^ (mul_22_8_n_967 ^ mul_22_8_n_968));
 assign mul_22_8_n_930 = ((mul_22_8_n_964 & mul_22_8_n_965) | (mul_22_8_n_963 & (mul_22_8_n_964 ^ mul_22_8_n_965)));
 assign mul_22_8_n_953 = (mul_22_8_n_963 ^ (mul_22_8_n_964 ^ mul_22_8_n_965));
 assign mul_22_8_n_929 = ((mul_22_8_n_961 & mul_22_8_n_962) | (mul_22_8_n_960 & (mul_22_8_n_961 ^ mul_22_8_n_962)));
 assign mul_22_8_n_954 = (mul_22_8_n_960 ^ (mul_22_8_n_961 ^ mul_22_8_n_962));
 assign mul_22_8_n_926 = ((mul_22_8_n_958 & mul_22_8_n_959) | (mul_22_8_n_957 & (mul_22_8_n_958 ^ mul_22_8_n_959)));
 assign mul_22_8_n_950 = (mul_22_8_n_957 ^ (mul_22_8_n_958 ^ mul_22_8_n_959));
 assign mul_22_8_n_925 = ((mul_22_8_n_955 & mul_22_8_n_956) | (mul_22_8_n_954 & (mul_22_8_n_955 ^ mul_22_8_n_956)));
 assign mul_22_8_n_949 = (mul_22_8_n_954 ^ (mul_22_8_n_955 ^ mul_22_8_n_956));
 assign mul_22_8_n_922 = ((mul_22_8_n_952 & mul_22_8_n_953) | (mul_22_8_n_951 & (mul_22_8_n_952 ^ mul_22_8_n_953)));
 assign mul_22_8_n_947 = (mul_22_8_n_951 ^ (mul_22_8_n_952 ^ mul_22_8_n_953));
 assign mul_22_8_n_919 = ((mul_22_8_n_949 & mul_22_8_n_950) | (mul_22_8_n_948 & (mul_22_8_n_949 ^ mul_22_8_n_950)));
 assign mul_22_8_n_946 = (mul_22_8_n_948 ^ (mul_22_8_n_949 ^ mul_22_8_n_950));
 assign mul_22_8_n_1316 = ((n_24 & n_52) | (n_54 & (n_24 ^ n_52)));
 assign mul_22_8_n_1291 = (n_54 ^ (n_24 ^ n_52));
 assign asc001_22_ = (mul_22_8_n_855 ^ mul_22_8_n_882);
 assign asc001_31_ = ~(mul_22_8_n_889 ^ mul_22_8_n_908);
 assign mul_22_8_n_908 = ((mul_22_8_n_1291 & n_154) | (mul_22_8_n_1315 & (mul_22_8_n_1291 ^ n_154)));
 assign asc001_30_ = (mul_22_8_n_1315 ^ (mul_22_8_n_1291 ^ n_154));
 assign asc001_29_ = ~(mul_22_8_n_893 ^ mul_22_8_n_904);
 assign asc001_27_ = ~(mul_22_8_n_875 ^ mul_22_8_n_903);
 assign mul_22_8_n_904 = (mul_22_8_n_898 & mul_22_8_n_886);
 assign mul_22_8_n_903 = ~(mul_22_8_n_838 | (mul_22_8_n_897 & mul_22_8_n_840));
 assign asc001_28_ = ~(mul_22_8_n_894 ^ mul_22_8_n_892);
 assign asc001_26_ = ~(mul_22_8_n_858 ^ mul_22_8_n_897);
 assign asc001_25_ = ~(mul_22_8_n_857 ^ mul_22_8_n_895);
 assign asc001_23_ = ~(mul_22_8_n_6 ^ mul_22_8_n_888);
 assign mul_22_8_n_898 = ~(~mul_22_8_n_892 & mul_22_8_n_884);
 assign mul_22_8_n_895 = ~(mul_22_8_n_834 | (mul_22_8_n_880 & mul_22_8_n_832));
 assign mul_22_8_n_894 = (mul_22_8_n_884 & mul_22_8_n_886);
 assign mul_22_8_n_893 = ~(~mul_22_8_n_887 | mul_22_8_n_885);
 assign mul_22_8_n_897 = ~(mul_22_8_n_861 & (mul_22_8_n_879 | mul_22_8_n_851));
 assign asc001_24_ = ~((mul_22_8_n_880 & ~mul_22_8_n_856) | (mul_22_8_n_879 & mul_22_8_n_856));
 assign asc001_21_ = ~(mul_22_8_n_854 ^ mul_22_8_n_881);
 assign mul_22_8_n_889 = ~(mul_22_8_n_1316 ^ mul_22_8_n_1292);
 assign mul_22_8_n_888 = ~(mul_22_8_n_835 & (mul_22_8_n_882 | mul_22_8_n_843));
 assign mul_22_8_n_892 = (mul_22_8_n_877 & (mul_22_8_n_883 & (mul_22_8_n_861 | mul_22_8_n_872)));
 assign mul_22_8_n_887 = ~(mul_22_8_n_1290 & mul_22_8_n_1314);
 assign mul_22_8_n_886 = ~(mul_22_8_n_1289 & mul_22_8_n_1313);
 assign mul_22_8_n_885 = ~(mul_22_8_n_1290 | mul_22_8_n_1314);
 assign mul_22_8_n_884 = (mul_22_8_n_1289 | mul_22_8_n_1313);
 assign mul_22_8_n_883 = ~(mul_22_8_n_880 & (~mul_22_8_n_872 & ~mul_22_8_n_851));
 assign mul_22_8_n_882 = ~(mul_22_8_n_862 | (mul_22_8_n_874 & mul_22_8_n_850));
 assign mul_22_8_n_881 = (~mul_22_8_n_842 | (mul_22_8_n_874 & mul_22_8_n_4));
 assign mul_22_8_n_879 = ~mul_22_8_n_880;
 assign mul_22_8_n_880 = ~(mul_22_8_n_873 & (mul_22_8_n_871 & (mul_22_8_n_863 | mul_22_8_n_864)));
 assign asc001_20_ = ~(mul_22_8_n_853 ^ mul_22_8_n_874);
 assign mul_22_8_n_877 = ~(mul_22_8_n_869 | (mul_22_8_n_870 & mul_22_8_n_838));
 assign asc001_19_ = ~(mul_22_8_n_5 ^ mul_22_8_n_868);
 assign mul_22_8_n_875 = ~(mul_22_8_n_869 | ~mul_22_8_n_870);
 assign mul_22_8_n_874 = ~(mul_22_8_n_863 & mul_22_8_n_867);
 assign mul_22_8_n_873 = (mul_22_8_n_867 | mul_22_8_n_864);
 assign mul_22_8_n_872 = ~(mul_22_8_n_870 & mul_22_8_n_840);
 assign mul_22_8_n_871 = ~(mul_22_8_n_848 | (mul_22_8_n_837 | (mul_22_8_n_862 & mul_22_8_n_859)));
 assign mul_22_8_n_870 = ~(mul_22_8_n_860 & n_75);
 assign mul_22_8_n_869 = ~(mul_22_8_n_860 | n_75);
 assign mul_22_8_n_868 = ~(n_49 & (mul_22_8_n_849 | n_48));
 assign mul_22_8_n_867 = ~(mul_22_8_n_847 | (n_38 | (mul_22_8_n_811 & mul_22_8_n_852)));
 assign asc001_18_ = (mul_22_8_n_819 ^ mul_22_8_n_849);
 assign asc001_17_ = ~(mul_22_8_n_807 ^ mul_22_8_n_846);
 assign mul_22_8_n_864 = ~(mul_22_8_n_859 & mul_22_8_n_850);
 assign mul_22_8_n_863 = ~(mul_22_8_n_836 & mul_22_8_n_852);
 assign mul_22_8_n_862 = ~(mul_22_8_n_844 & (mul_22_8_n_841 | mul_22_8_n_842));
 assign mul_22_8_n_861 = ~(mul_22_8_n_845 | (mul_22_8_n_833 & mul_22_8_n_834));
 assign mul_22_8_n_860 = ~mul_22_8_n_1288;
 assign mul_22_8_n_858 = ~(~mul_22_8_n_838 & mul_22_8_n_840);
 assign mul_22_8_n_857 = ~(mul_22_8_n_845 | ~mul_22_8_n_833);
 assign mul_22_8_n_856 = ~(~mul_22_8_n_834 & mul_22_8_n_832);
 assign mul_22_8_n_859 = ~(mul_22_8_n_839 | mul_22_8_n_843);
 assign mul_22_8_n_855 = ~(~mul_22_8_n_843 & mul_22_8_n_835);
 assign mul_22_8_n_854 = ~(mul_22_8_n_844 & ~mul_22_8_n_841);
 assign mul_22_8_n_853 = ~(mul_22_8_n_4 & mul_22_8_n_842);
 assign mul_22_8_n_848 = ~(mul_22_8_n_839 | mul_22_8_n_835);
 assign mul_22_8_n_847 = ~(n_28 | n_49);
 assign mul_22_8_n_852 = ~(n_28 | n_48);
 assign mul_22_8_n_851 = ~(mul_22_8_n_833 & mul_22_8_n_832);
 assign mul_22_8_n_846 = ~(n_45 & (mul_22_8_n_827 | n_46));
 assign mul_22_8_n_850 = ~(~mul_22_8_n_4 | mul_22_8_n_841);
 assign mul_22_8_n_849 = ~(mul_22_8_n_836 | mul_22_8_n_811);
 assign mul_22_8_n_845 = ~(mul_22_8_n_824 | n_78);
 assign mul_22_8_n_844 = ~(mul_22_8_n_1282 & n_37);
 assign mul_22_8_n_843 = ~(n_72 | mul_22_8_n_1307);
 assign mul_22_8_n_842 = ~(n_36 & n_81);
 assign mul_22_8_n_841 = ~(mul_22_8_n_1282 | n_37);
 assign mul_22_8_n_840 = ~(mul_22_8_n_828 & mul_22_8_n_829);
 assign mul_22_8_n_839 = ~(mul_22_8_n_1284 | n_73);
 assign mul_22_8_n_838 = ~(mul_22_8_n_828 | mul_22_8_n_829);
 assign asc001_15_ = ~(mul_22_8_n_806 ^ mul_22_8_n_821);
 assign mul_22_8_n_837 = (mul_22_8_n_1284 & n_73);
 assign mul_22_8_n_836 = ~(n_31 | (n_46 | mul_22_8_n_827));
 assign mul_22_8_n_835 = ~(n_72 & mul_22_8_n_1307);
 assign mul_22_8_n_834 = ~(mul_22_8_n_823 | mul_22_8_n_826);
 assign mul_22_8_n_833 = ~(mul_22_8_n_824 & n_78);
 assign mul_22_8_n_832 = ~(mul_22_8_n_823 & mul_22_8_n_826);
 assign mul_22_8_n_831 = ~(mul_22_8_n_1280 | mul_22_8_n_1304);
 assign mul_22_8_n_829 = ~mul_22_8_n_1311;
 assign mul_22_8_n_827 = ~(mul_22_8_n_817 | (mul_22_8_n_818 | (n_27 & mul_22_8_n_812)));
 assign mul_22_8_n_826 = ~mul_22_8_n_1309;
 assign mul_22_8_n_825 = ~mul_22_8_n_1310;
 assign mul_22_8_n_824 = ~mul_22_8_n_1286;
 assign mul_22_8_n_822 = ~mul_22_8_n_1312;
 assign mul_22_8_n_821 = ~(n_26 | (mul_22_8_n_814 & n_42));
 assign asc001_14_ = ~(mul_22_8_n_803 ^ mul_22_8_n_814);
 assign mul_22_8_n_819 = ~(n_49 & ~n_48);
 assign mul_22_8_n_818 = ~(mul_22_8_n_804 & (n_60 & (mul_22_8_n_810 | mul_22_8_n_805)));
 assign mul_22_8_n_817 = (n_66 & mul_22_8_n_812);
 assign mul_22_8_n_816 = ~(mul_22_8_n_1279 & mul_22_8_n_1303);
 assign mul_22_8_n_815 = ~(mul_22_8_n_1279 | mul_22_8_n_1303);
 assign mul_22_8_n_814 = ~(mul_22_8_n_810 & (mul_22_8_n_785 | mul_22_8_n_809));
 assign asc001_13_ = ~(mul_22_8_n_802 ^ mul_22_8_n_789);
 assign mul_22_8_n_812 = ~(mul_22_8_n_805 | mul_22_8_n_809);
 assign mul_22_8_n_811 = ~(n_61 & (n_31 | n_45));
 assign mul_22_8_n_810 = ~(n_47 | (n_62 & n_34));
 assign mul_22_8_n_808 = ~(~n_46 & n_45);
 assign mul_22_8_n_807 = ~(~n_31 & n_61);
 assign mul_22_8_n_809 = ~(n_62 & n_63);
 assign mul_22_8_n_806 = (n_50 & n_60);
 assign mul_22_8_n_804 = ~(n_50 & n_26);
 assign mul_22_8_n_805 = ~(n_50 & n_42);
 assign mul_22_8_n_803 = ~(n_42 & ~n_26);
 assign mul_22_8_n_802 = ~(n_47 | ~n_62);
 assign mul_22_8_n_801 = ~(mul_22_8_n_1278 & mul_22_8_n_1302);
 assign mul_22_8_n_800 = ~(mul_22_8_n_1276 & mul_22_8_n_1300);
 assign mul_22_8_n_799 = ~(mul_22_8_n_1277 & mul_22_8_n_1301);
 assign mul_22_8_n_798 = ~(mul_22_8_n_1278 | mul_22_8_n_1302);
 assign mul_22_8_n_797 = ~(mul_22_8_n_1277 | mul_22_8_n_1301);
 assign mul_22_8_n_796 = ~(mul_22_8_n_787 | mul_22_8_n_788);
 assign mul_22_8_n_795 = ~(mul_22_8_n_786 & mul_22_8_n_774);
 assign asc001_11_ = (n_64 ^ mul_22_8_n_1);
 assign asc001_12_ = ~(mul_22_8_n_783 ^ mul_22_8_n_785);
 assign mul_22_8_n_794 = ~(mul_22_8_n_786 | mul_22_8_n_774);
 assign mul_22_8_n_789 = ~(n_34 | (~mul_22_8_n_785 & n_63));
 assign mul_22_8_n_793 = (mul_22_8_n_1276 | mul_22_8_n_1300);
 assign mul_22_8_n_792 = ~(mul_22_8_n_787 & mul_22_8_n_788);
 assign mul_22_8_n_788 = ~mul_22_8_n_1299;
 assign mul_22_8_n_787 = ~mul_22_8_n_1275;
 assign mul_22_8_n_786 = ~mul_22_8_n_1274;
 assign mul_22_8_n_785 = ~(n_27 | n_66);
 assign asc001_10_ = (mul_22_8_n_770 ^ n_86);
 assign mul_22_8_n_783 = ~(n_34 | ~n_63);
 assign mul_22_8_n_782 = ~(mul_22_8_n_771 & (mul_22_8_n_767 & (mul_22_8_n_776 | mul_22_8_n_772)));
 assign mul_22_8_n_781 = ~(mul_22_8_n_775 | mul_22_8_n_760);
 assign mul_22_8_n_780 = ~(mul_22_8_n_775 & mul_22_8_n_760);
 assign mul_22_8_n_779 = ~(mul_22_8_n_773 & mul_22_8_n_776);
 assign asc001_9_ = ~(mul_22_8_n_768 ^ mul_22_8_n_757);
 assign mul_22_8_n_775 = ~mul_22_8_n_1273;
 assign mul_22_8_n_777 = ~(mul_22_8_n_773 | mul_22_8_n_772);
 assign mul_22_8_n_776 = ~(mul_22_8_n_762 | (mul_22_8_n_761 & mul_22_8_n_752));
 assign mul_22_8_n_774 = ~mul_22_8_n_1298;
 assign mul_22_8_n_771 = ~(~mul_22_8_n_766 & mul_22_8_n_765);
 assign mul_22_8_n_773 = ~(mul_22_8_n_756 & mul_22_8_n_761);
 assign mul_22_8_n_772 = (mul_22_8_n_764 | mul_22_8_n_763);
 assign mul_22_8_n_770 = ~(n_67 | ~n_65);
 assign mul_22_8_n_769 = (mul_22_8_n_765 & mul_22_8_n_767);
 assign mul_22_8_n_768 = ~(mul_22_8_n_762 | ~mul_22_8_n_761);
 assign mul_22_8_n_767 = ~(mul_22_8_n_1272 & mul_22_8_n_1296);
 assign mul_22_8_n_766 = ~(mul_22_8_n_1271 & mul_22_8_n_1295);
 assign mul_22_8_n_765 = ~mul_22_8_n_764;
 assign mul_22_8_n_764 = ~(mul_22_8_n_1272 | mul_22_8_n_1296);
 assign mul_22_8_n_763 = ~(mul_22_8_n_1271 | mul_22_8_n_1295);
 assign mul_22_8_n_762 = ~(mul_22_8_n_759 | mul_22_8_n_749);
 assign mul_22_8_n_761 = ~(mul_22_8_n_759 & mul_22_8_n_749);
 assign mul_22_8_n_760 = ~mul_22_8_n_1297;
 assign mul_22_8_n_759 = ~mul_22_8_n_1270;
 assign asc001_8_ = ~(mul_22_8_n_755 ^ mul_22_8_n_754);
 assign mul_22_8_n_757 = ~(mul_22_8_n_756 | mul_22_8_n_752);
 assign mul_22_8_n_756 = ~(mul_22_8_n_754 | mul_22_8_n_751);
 assign mul_22_8_n_755 = ~(mul_22_8_n_751 | mul_22_8_n_752);
 assign mul_22_8_n_754 = ~(mul_22_8_n_748 | (mul_22_8_n_747 | (mul_22_8_n_734 & mul_22_8_n_744)));
 assign asc001_7_ = ~(mul_22_8_n_743 ^ mul_22_8_n_746);
 assign mul_22_8_n_752 = ~(mul_22_8_n_745 | mul_22_8_n_735);
 assign mul_22_8_n_751 = (mul_22_8_n_745 & mul_22_8_n_735);
 assign asc001_6_ = ~(mul_22_8_n_737 ^ mul_22_8_n_742);
 assign mul_22_8_n_749 = ~mul_22_8_n_1294;
 assign mul_22_8_n_748 = ~(mul_22_8_n_741 & (mul_22_8_n_739 | mul_22_8_n_740));
 assign mul_22_8_n_747 = (mul_22_8_n_733 & mul_22_8_n_744);
 assign mul_22_8_n_746 = ~(mul_22_8_n_740 & (mul_22_8_n_737 | mul_22_8_n_738));
 assign mul_22_8_n_745 = ~mul_22_8_n_911;
 assign mul_22_8_n_744 = ~(mul_22_8_n_739 | mul_22_8_n_738);
 assign mul_22_8_n_743 = ~(~mul_22_8_n_739 & mul_22_8_n_741);
 assign mul_22_8_n_742 = ~(mul_22_8_n_738 | ~mul_22_8_n_740);
 assign mul_22_8_n_741 = ~(mul_22_8_n_912 & mul_22_8_n_915);
 assign mul_22_8_n_740 = ~(mul_22_8_n_914 & mul_22_8_n_1293);
 assign mul_22_8_n_739 = ~(mul_22_8_n_912 | mul_22_8_n_915);
 assign mul_22_8_n_738 = ~(mul_22_8_n_914 | mul_22_8_n_1293);
 assign asc001_5_ = ~(mul_22_8_n_728 ^ mul_22_8_n_732);
 assign mul_22_8_n_737 = ~(mul_22_8_n_733 | mul_22_8_n_734);
 assign mul_22_8_n_735 = ~mul_22_8_n_913;
 assign mul_22_8_n_734 = ~(mul_22_8_n_731 & (mul_22_8_n_725 | mul_22_8_n_730));
 assign mul_22_8_n_733 = ~(mul_22_8_n_726 | mul_22_8_n_730);
 assign mul_22_8_n_732 = ~(mul_22_8_n_730 | ~mul_22_8_n_731);
 assign mul_22_8_n_731 = ~(mul_22_8_n_916 & mul_22_8_n_918);
 assign mul_22_8_n_730 = ~(mul_22_8_n_916 | mul_22_8_n_918);
 assign asc001_4_ = ~(mul_22_8_n_723 ^ mul_22_8_n_727);
 assign mul_22_8_n_728 = (mul_22_8_n_726 & mul_22_8_n_725);
 assign mul_22_8_n_727 = ~(mul_22_8_n_725 & mul_22_8_n_724);
 assign mul_22_8_n_726 = ~(mul_22_8_n_723 & mul_22_8_n_724);
 assign mul_22_8_n_725 = ~(mul_22_8_n_691 & mul_22_8_n_917);
 assign mul_22_8_n_724 = (mul_22_8_n_691 | mul_22_8_n_917);
 assign asc001_3_ = ~(mul_22_8_n_719 ^ mul_22_8_n_720);
 assign mul_22_8_n_723 = ~(mul_22_8_n_721 & (mul_22_8_n_718 & (mul_22_8_n_717 | mul_22_8_n_715)));
 assign mul_22_8_n_721 = ~(mul_22_8_n_673 & ~mul_22_8_n_717);
 assign mul_22_8_n_720 = ~(mul_22_8_n_718 & ~mul_22_8_n_717);
 assign mul_22_8_n_719 = ~(~mul_22_8_n_673 & mul_22_8_n_715);
 assign mul_22_8_n_718 = ~(mul_22_8_n_714 & mul_22_8_n_683);
 assign mul_22_8_n_717 = ~(mul_22_8_n_714 | mul_22_8_n_683);
 assign asc001_2_ = ~(mul_22_8_n_665 ^ mul_22_8_n_684);
 assign mul_22_8_n_715 = ~(mul_22_8_n_682 & mul_22_8_n_665);
 assign mul_22_8_n_713 = ~(mul_22_8_n_675 ^ mul_22_8_n_671);
 assign mul_22_8_n_712 = ~(mul_22_8_n_672 ^ mul_22_8_n_558);
 assign mul_22_8_n_711 = (mul_22_8_n_681 ^ mul_22_8_n_559);
 assign mul_22_8_n_710 = (mul_22_8_n_669 ^ mul_22_8_n_560);
 assign mul_22_8_n_709 = (mul_22_8_n_561 ^ mul_22_8_n_680);
 assign mul_22_8_n_708 = (mul_22_8_n_670 ^ mul_22_8_n_562);
 assign mul_22_8_n_714 = (mul_22_8_n_667 ^ mul_22_8_n_413);
 assign mul_22_8_n_707 = (mul_22_8_n_563 ^ mul_22_8_n_418);
 assign mul_22_8_n_706 = (mul_22_8_n_666 ^ mul_22_8_n_439);
 assign mul_22_8_n_705 = (mul_22_8_n_411 ^ mul_22_8_n_668);
 assign mul_22_8_n_704 = (mul_22_8_n_674 ^ mul_22_8_n_412);
 assign mul_22_8_n_703 = (mul_22_8_n_679 ^ mul_22_8_n_438);
 assign mul_22_8_n_702 = (mul_22_8_n_676 ^ mul_22_8_n_415);
 assign mul_22_8_n_701 = (mul_22_8_n_678 ^ mul_22_8_n_416);
 assign mul_22_8_n_700 = (mul_22_8_n_677 ^ mul_22_8_n_414);
 assign mul_22_8_n_699 = ~(mul_22_8_n_438 | mul_22_8_n_679);
 assign mul_22_8_n_698 = ~(mul_22_8_n_415 | mul_22_8_n_676);
 assign mul_22_8_n_697 = ~(mul_22_8_n_414 | mul_22_8_n_677);
 assign mul_22_8_n_696 = ~(mul_22_8_n_416 | mul_22_8_n_678);
 assign mul_22_8_n_695 = ~(mul_22_8_n_411 | mul_22_8_n_668);
 assign mul_22_8_n_694 = ~(mul_22_8_n_412 | mul_22_8_n_674);
 assign mul_22_8_n_693 = ~(mul_22_8_n_560 | mul_22_8_n_669);
 assign mul_22_8_n_692 = ~(mul_22_8_n_439 | mul_22_8_n_666);
 assign mul_22_8_n_690 = ~(mul_22_8_n_675 | ~mul_22_8_n_671);
 assign mul_22_8_n_689 = ~(mul_22_8_n_562 | mul_22_8_n_670);
 assign mul_22_8_n_688 = ~(mul_22_8_n_672 | ~mul_22_8_n_558);
 assign asc001_1_ = ~(mul_22_8_n_665 | (mul_22_8_n_440 & mul_22_8_n_360));
 assign mul_22_8_n_686 = ~(mul_22_8_n_559 | mul_22_8_n_681);
 assign mul_22_8_n_685 = ~(mul_22_8_n_561 | mul_22_8_n_680);
 assign mul_22_8_n_691 = ~(mul_22_8_n_413 | mul_22_8_n_667);
 assign mul_22_8_n_684 = ~(mul_22_8_n_682 & ~mul_22_8_n_673);
 assign mul_22_8_n_664 = ~((mul_22_8_n_235 | mul_22_8_n_251) & (mul_22_8_n_369 | mul_22_8_n_250));
 assign mul_22_8_n_663 = ~((mul_22_8_n_232 | mul_22_8_n_323) & (mul_22_8_n_366 | mul_22_8_n_320));
 assign mul_22_8_n_662 = ~((mul_22_8_n_238 | mul_22_8_n_126) & (mul_22_8_n_372 | mul_22_8_n_115));
 assign mul_22_8_n_661 = ~((n_155 | mul_22_8_n_122) & (mul_22_8_n_377 | mul_22_8_n_129));
 assign mul_22_8_n_660 = ~((mul_22_8_n_237 | mul_22_8_n_186) & (mul_22_8_n_371 | mul_22_8_n_185));
 assign mul_22_8_n_659 = ~((mul_22_8_n_234 | mul_22_8_n_355) & (mul_22_8_n_368 | mul_22_8_n_325));
 assign mul_22_8_n_658 = ~((mul_22_8_n_233 | mul_22_8_n_137) & (mul_22_8_n_367 | mul_22_8_n_128));
 assign mul_22_8_n_657 = ~((mul_22_8_n_236 | mul_22_8_n_199) & (mul_22_8_n_370 | mul_22_8_n_198));
 assign mul_22_8_n_656 = ~((mul_22_8_n_236 | mul_22_8_n_304) & (mul_22_8_n_370 | mul_22_8_n_286));
 assign mul_22_8_n_655 = ~((mul_22_8_n_232 | mul_22_8_n_318) & (mul_22_8_n_366 | mul_22_8_n_323));
 assign mul_22_8_n_654 = ~((mul_22_8_n_242 | mul_22_8_n_81) & (mul_22_8_n_376 | mul_22_8_n_82));
 assign mul_22_8_n_653 = ~((mul_22_8_n_232 | mul_22_8_n_264) & (mul_22_8_n_366 | mul_22_8_n_246));
 assign mul_22_8_n_652 = ~((mul_22_8_n_244 | mul_22_8_n_254) & (mul_22_8_n_379 | mul_22_8_n_263));
 assign mul_22_8_n_651 = ~((mul_22_8_n_232 | mul_22_8_n_246) & (mul_22_8_n_366 | mul_22_8_n_262));
 assign mul_22_8_n_650 = ~((mul_22_8_n_237 | mul_22_8_n_300) & (mul_22_8_n_371 | mul_22_8_n_281));
 assign mul_22_8_n_649 = ~((n_155 | mul_22_8_n_98) & (mul_22_8_n_377 | mul_22_8_n_110));
 assign mul_22_8_n_648 = ~((mul_22_8_n_236 | mul_22_8_n_319) & (mul_22_8_n_370 | mul_22_8_n_303));
 assign mul_22_8_n_647 = ~((mul_22_8_n_241 | mul_22_8_n_114) & (mul_22_8_n_375 | mul_22_8_n_113));
 assign mul_22_8_n_646 = ~(mul_22_8_n_364 & (mul_22_8_n_245 | (mul_22_8_n_51 | mul_22_8_n_226)));
 assign mul_22_8_n_645 = ~((mul_22_8_n_232 | mul_22_8_n_229) & (mul_22_8_n_366 | mul_22_8_n_318));
 assign mul_22_8_n_644 = ~((mul_22_8_n_233 | mul_22_8_n_225) & (mul_22_8_n_367 | mul_22_8_n_301));
 assign mul_22_8_n_643 = ~((mul_22_8_n_234 | mul_22_8_n_223) & (mul_22_8_n_368 | mul_22_8_n_350));
 assign mul_22_8_n_642 = ~((mul_22_8_n_235 | mul_22_8_n_222) & (mul_22_8_n_369 | mul_22_8_n_348));
 assign mul_22_8_n_641 = ~((mul_22_8_n_236 | mul_22_8_n_214) & (mul_22_8_n_370 | mul_22_8_n_319));
 assign mul_22_8_n_640 = ~((mul_22_8_n_244 | mul_22_8_n_263) & (mul_22_8_n_379 | mul_22_8_n_210));
 assign mul_22_8_n_639 = ~((mul_22_8_n_237 | mul_22_8_n_209) & (mul_22_8_n_371 | mul_22_8_n_300));
 assign mul_22_8_n_638 = ~((mul_22_8_n_238 | mul_22_8_n_208) & (mul_22_8_n_372 | mul_22_8_n_275));
 assign mul_22_8_n_637 = ~((mul_22_8_n_0 | mul_22_8_n_194) & (mul_22_8_n_378 | mul_22_8_n_207));
 assign mul_22_8_n_636 = ~((mul_22_8_n_244 | mul_22_8_n_206) & (mul_22_8_n_379 | mul_22_8_n_254));
 assign mul_22_8_n_635 = ~((mul_22_8_n_239 | mul_22_8_n_213) & (mul_22_8_n_373 | mul_22_8_n_324));
 assign mul_22_8_n_634 = ~((n_155 | mul_22_8_n_129) & (mul_22_8_n_377 | mul_22_8_n_230));
 assign mul_22_8_n_633 = ~((mul_22_8_n_240 | mul_22_8_n_60) & (mul_22_8_n_374 | mul_22_8_n_190));
 assign mul_22_8_n_632 = ~((mul_22_8_n_242 | mul_22_8_n_100) & (mul_22_8_n_376 | mul_22_8_n_68));
 assign mul_22_8_n_631 = ~((mul_22_8_n_0 | mul_22_8_n_67) & (mul_22_8_n_378 | mul_22_8_n_166));
 assign mul_22_8_n_630 = ~((mul_22_8_n_241 | mul_22_8_n_77) & (mul_22_8_n_375 | mul_22_8_n_66));
 assign mul_22_8_n_629 = ~((mul_22_8_n_241 | mul_22_8_n_64) & (mul_22_8_n_375 | mul_22_8_n_138));
 assign mul_22_8_n_628 = ~((mul_22_8_n_240 | mul_22_8_n_85) & (mul_22_8_n_374 | mul_22_8_n_63));
 assign mul_22_8_n_627 = ~((mul_22_8_n_239 | mul_22_8_n_95) & (mul_22_8_n_373 | mul_22_8_n_62));
 assign mul_22_8_n_626 = ~((mul_22_8_n_238 | mul_22_8_n_108) & (mul_22_8_n_372 | mul_22_8_n_61));
 assign mul_22_8_n_625 = ~((n_155 | mul_22_8_n_69) & (mul_22_8_n_377 | mul_22_8_n_98));
 assign mul_22_8_n_624 = ~((mul_22_8_n_242 | mul_22_8_n_59) & (mul_22_8_n_376 | mul_22_8_n_97));
 assign mul_22_8_n_623 = ~((mul_22_8_n_237 | mul_22_8_n_112) & (mul_22_8_n_371 | mul_22_8_n_58));
 assign mul_22_8_n_622 = ~((mul_22_8_n_236 | mul_22_8_n_123) & (mul_22_8_n_370 | mul_22_8_n_57));
 assign mul_22_8_n_621 = ~((mul_22_8_n_235 | mul_22_8_n_130) & (mul_22_8_n_369 | mul_22_8_n_56));
 assign mul_22_8_n_620 = ~((mul_22_8_n_234 | mul_22_8_n_139) & (mul_22_8_n_368 | mul_22_8_n_54));
 assign mul_22_8_n_619 = ~((mul_22_8_n_234 | mul_22_8_n_155) & (mul_22_8_n_368 | mul_22_8_n_154));
 assign mul_22_8_n_618 = ~((mul_22_8_n_233 | mul_22_8_n_147) & (mul_22_8_n_367 | mul_22_8_n_52));
 assign mul_22_8_n_617 = ~((mul_22_8_n_239 | mul_22_8_n_324) & (mul_22_8_n_373 | mul_22_8_n_76));
 assign mul_22_8_n_616 = ~((mul_22_8_n_232 | mul_22_8_n_262) & (mul_22_8_n_366 | mul_22_8_n_165));
 assign mul_22_8_n_615 = ~((mul_22_8_n_234 | mul_22_8_n_350) & (mul_22_8_n_368 | mul_22_8_n_354));
 assign mul_22_8_n_614 = ~((mul_22_8_n_238 | mul_22_8_n_127) & (mul_22_8_n_372 | mul_22_8_n_126));
 assign mul_22_8_n_613 = ~((mul_22_8_n_235 | mul_22_8_n_348) & (mul_22_8_n_369 | mul_22_8_n_321));
 assign mul_22_8_n_612 = ~((mul_22_8_n_239 | mul_22_8_n_106) & (mul_22_8_n_373 | mul_22_8_n_107));
 assign mul_22_8_n_611 = ~((mul_22_8_n_234 | mul_22_8_n_193) & (mul_22_8_n_368 | mul_22_8_n_172));
 assign mul_22_8_n_610 = ~((mul_22_8_n_232 | mul_22_8_n_320) & (mul_22_8_n_366 | mul_22_8_n_302));
 assign mul_22_8_n_609 = ~((mul_22_8_n_232 | mul_22_8_n_296) & (mul_22_8_n_366 | mul_22_8_n_295));
 assign mul_22_8_n_608 = ~((mul_22_8_n_239 | mul_22_8_n_78) & (mul_22_8_n_373 | mul_22_8_n_182));
 assign mul_22_8_n_607 = ~((mul_22_8_n_240 | mul_22_8_n_157) & (mul_22_8_n_374 | mul_22_8_n_133));
 assign mul_22_8_n_606 = ~((mul_22_8_n_241 | mul_22_8_n_113) & (mul_22_8_n_375 | mul_22_8_n_102));
 assign mul_22_8_n_605 = ~((mul_22_8_n_235 | mul_22_8_n_164) & (mul_22_8_n_369 | mul_22_8_n_143));
 assign mul_22_8_n_604 = ~((mul_22_8_n_235 | mul_22_8_n_250) & (mul_22_8_n_369 | mul_22_8_n_343));
 assign mul_22_8_n_603 = ~((mul_22_8_n_235 | mul_22_8_n_289) & (mul_22_8_n_369 | mul_22_8_n_271));
 assign mul_22_8_n_602 = ~((mul_22_8_n_242 | mul_22_8_n_83) & (mul_22_8_n_376 | mul_22_8_n_81));
 assign mul_22_8_n_601 = ~((n_155 | mul_22_8_n_109) & (mul_22_8_n_377 | mul_22_8_n_121));
 assign mul_22_8_n_600 = ~((mul_22_8_n_233 | mul_22_8_n_278) & (mul_22_8_n_367 | mul_22_8_n_277));
 assign mul_22_8_n_599 = ~((mul_22_8_n_236 | mul_22_8_n_136) & (mul_22_8_n_370 | mul_22_8_n_123));
 assign mul_22_8_n_598 = ~((mul_22_8_n_233 | mul_22_8_n_276) & (mul_22_8_n_367 | mul_22_8_n_359));
 assign mul_22_8_n_597 = ~((mul_22_8_n_0 | mul_22_8_n_178) & (mul_22_8_n_378 | mul_22_8_n_194));
 assign mul_22_8_n_596 = ~((mul_22_8_n_237 | mul_22_8_n_160) & (mul_22_8_n_371 | mul_22_8_n_159));
 assign mul_22_8_n_595 = ~((mul_22_8_n_237 | mul_22_8_n_282) & (mul_22_8_n_371 | mul_22_8_n_258));
 assign mul_22_8_n_594 = ~((mul_22_8_n_239 | mul_22_8_n_151) & (mul_22_8_n_373 | mul_22_8_n_132));
 assign mul_22_8_n_593 = ~((mul_22_8_n_234 | mul_22_8_n_256) & (mul_22_8_n_368 | mul_22_8_n_344));
 assign mul_22_8_n_592 = ~((mul_22_8_n_236 | mul_22_8_n_286) & (mul_22_8_n_370 | mul_22_8_n_287));
 assign mul_22_8_n_591 = ~((mul_22_8_n_234 | mul_22_8_n_96) & (mul_22_8_n_368 | mul_22_8_n_192));
 assign mul_22_8_n_590 = ~((mul_22_8_n_234 | mul_22_8_n_192) & (mul_22_8_n_368 | mul_22_8_n_193));
 assign mul_22_8_n_589 = ~((mul_22_8_n_233 | mul_22_8_n_359) & (mul_22_8_n_367 | mul_22_8_n_270));
 assign mul_22_8_n_588 = ~((mul_22_8_n_238 | mul_22_8_n_201) & (mul_22_8_n_372 | mul_22_8_n_169));
 assign mul_22_8_n_587 = ~((n_155 | mul_22_8_n_121) & (mul_22_8_n_377 | mul_22_8_n_122));
 assign mul_22_8_n_586 = ~((mul_22_8_n_238 | mul_22_8_n_253) & (mul_22_8_n_372 | mul_22_8_n_140));
 assign mul_22_8_n_585 = ~((mul_22_8_n_240 | mul_22_8_n_94) & (mul_22_8_n_374 | mul_22_8_n_85));
 assign mul_22_8_n_584 = ~((mul_22_8_n_235 | mul_22_8_n_343) & (mul_22_8_n_369 | mul_22_8_n_148));
 assign mul_22_8_n_583 = ~((mul_22_8_n_235 | mul_22_8_n_321) & (mul_22_8_n_369 | mul_22_8_n_322));
 assign mul_22_8_n_582 = ~((mul_22_8_n_233 | mul_22_8_n_161) & (mul_22_8_n_367 | mul_22_8_n_162));
 assign mul_22_8_n_581 = ~((mul_22_8_n_236 | mul_22_8_n_303) & (mul_22_8_n_370 | mul_22_8_n_304));
 assign mul_22_8_n_580 = ~((mul_22_8_n_232 | mul_22_8_n_279) & (mul_22_8_n_366 | mul_22_8_n_265));
 assign mul_22_8_n_579 = ~((mul_22_8_n_233 | mul_22_8_n_357) & (mul_22_8_n_367 | mul_22_8_n_276));
 assign mul_22_8_n_578 = ~((n_155 | mul_22_8_n_110) & (mul_22_8_n_377 | mul_22_8_n_109));
 assign mul_22_8_n_577 = ~((mul_22_8_n_242 | mul_22_8_n_97) & (mul_22_8_n_376 | mul_22_8_n_84));
 assign mul_22_8_n_576 = ~((mul_22_8_n_233 | mul_22_8_n_128) & (mul_22_8_n_367 | mul_22_8_n_202));
 assign mul_22_8_n_575 = ~((mul_22_8_n_0 | mul_22_8_n_177) & (mul_22_8_n_378 | mul_22_8_n_178));
 assign mul_22_8_n_574 = ~((mul_22_8_n_239 | mul_22_8_n_117) & (mul_22_8_n_373 | mul_22_8_n_106));
 assign mul_22_8_n_573 = ~((mul_22_8_n_232 | mul_22_8_n_313) & (mul_22_8_n_366 | mul_22_8_n_296));
 assign mul_22_8_n_572 = ~((mul_22_8_n_237 | mul_22_8_n_159) & (mul_22_8_n_371 | mul_22_8_n_142));
 assign mul_22_8_n_571 = ~((mul_22_8_n_233 | mul_22_8_n_203) & (mul_22_8_n_367 | mul_22_8_n_180));
 assign mul_22_8_n_570 = ~((mul_22_8_n_234 | mul_22_8_n_354) & (mul_22_8_n_368 | mul_22_8_n_355));
 assign mul_22_8_n_569 = ~((mul_22_8_n_236 | mul_22_8_n_111) & (mul_22_8_n_370 | mul_22_8_n_199));
 assign mul_22_8_n_568 = ~((mul_22_8_n_236 | mul_22_8_n_103) & (mul_22_8_n_370 | mul_22_8_n_111));
 assign mul_22_8_n_567 = ~((mul_22_8_n_236 | mul_22_8_n_135) & (mul_22_8_n_370 | mul_22_8_n_136));
 assign mul_22_8_n_566 = ~((mul_22_8_n_232 | mul_22_8_n_187) & (mul_22_8_n_366 | mul_22_8_n_188));
 assign mul_22_8_n_565 = ~((mul_22_8_n_238 | mul_22_8_n_275) & (mul_22_8_n_372 | mul_22_8_n_252));
 assign mul_22_8_n_564 = ~((mul_22_8_n_237 | mul_22_8_n_259) & (mul_22_8_n_371 | mul_22_8_n_339));
 assign mul_22_8_n_683 = ~((mul_22_8_n_232 | mul_22_8_n_152) & (mul_22_8_n_366 | mul_22_8_n_53));
 assign mul_22_8_n_563 = ~(mul_22_8_n_430 & {in2[31]});
 assign mul_22_8_n_682 = ~(mul_22_8_n_417 & mul_22_8_n_394);
 assign mul_22_8_n_681 = ~(mul_22_8_n_432 & {in2[9]});
 assign mul_22_8_n_680 = ~(mul_22_8_n_424 & {in2[11]});
 assign mul_22_8_n_679 = ~(mul_22_8_n_436 & {in2[13]});
 assign mul_22_8_n_678 = ~(mul_22_8_n_431 & {in2[15]});
 assign mul_22_8_n_677 = ~(mul_22_8_n_423 & {in2[17]});
 assign mul_22_8_n_676 = ~(mul_22_8_n_422 & {in2[19]});
 assign mul_22_8_n_675 = ~(mul_22_8_n_433 & {in2[21]});
 assign mul_22_8_n_674 = ~(mul_22_8_n_425 & {in2[7]});
 assign mul_22_8_n_673 = ~(mul_22_8_n_417 | mul_22_8_n_394);
 assign mul_22_8_n_672 = ~(mul_22_8_n_428 & {in2[23]});
 assign mul_22_8_n_671 = ~((mul_22_8_n_232 | mul_22_8_n_314) & (mul_22_8_n_366 | mul_22_8_n_313));
 assign mul_22_8_n_670 = ~(mul_22_8_n_434 & {in2[25]});
 assign mul_22_8_n_669 = ~(mul_22_8_n_426 & {in2[27]});
 assign mul_22_8_n_668 = ~(mul_22_8_n_429 & {in2[29]});
 assign mul_22_8_n_667 = ~(mul_22_8_n_427 & {in2[3]});
 assign mul_22_8_n_666 = ~(mul_22_8_n_435 & {in2[5]});
 assign mul_22_8_n_665 = ~(mul_22_8_n_440 | mul_22_8_n_360);
 assign mul_22_8_n_557 = ~((mul_22_8_n_233 | mul_22_8_n_162) & (mul_22_8_n_367 | mul_22_8_n_147));
 assign mul_22_8_n_556 = ~((mul_22_8_n_236 | mul_22_8_n_191) & (mul_22_8_n_370 | mul_22_8_n_135));
 assign mul_22_8_n_555 = ~((mul_22_8_n_232 | mul_22_8_n_329) & (mul_22_8_n_366 | mul_22_8_n_314));
 assign mul_22_8_n_554 = ~((mul_22_8_n_234 | mul_22_8_n_290) & (mul_22_8_n_368 | mul_22_8_n_273));
 assign mul_22_8_n_553 = ~((mul_22_8_n_237 | mul_22_8_n_124) & (mul_22_8_n_371 | mul_22_8_n_112));
 assign mul_22_8_n_552 = ~((mul_22_8_n_238 | mul_22_8_n_170) & (mul_22_8_n_372 | mul_22_8_n_145));
 assign mul_22_8_n_551 = ~((mul_22_8_n_234 | mul_22_8_n_154) & (mul_22_8_n_368 | mul_22_8_n_139));
 assign mul_22_8_n_550 = ~((mul_22_8_n_239 | mul_22_8_n_131) & (mul_22_8_n_373 | mul_22_8_n_118));
 assign mul_22_8_n_549 = ~((mul_22_8_n_235 | mul_22_8_n_272) & (mul_22_8_n_369 | mul_22_8_n_251));
 assign mul_22_8_n_548 = ~((mul_22_8_n_240 | mul_22_8_n_104) & (mul_22_8_n_374 | mul_22_8_n_93));
 assign mul_22_8_n_547 = ~((mul_22_8_n_241 | mul_22_8_n_80) & (mul_22_8_n_375 | mul_22_8_n_77));
 assign mul_22_8_n_546 = ~((mul_22_8_n_235 | mul_22_8_n_271) & (mul_22_8_n_369 | mul_22_8_n_272));
 assign mul_22_8_n_545 = ~((mul_22_8_n_233 | mul_22_8_n_312) & (mul_22_8_n_367 | mul_22_8_n_294));
 assign mul_22_8_n_544 = ~((mul_22_8_n_236 | mul_22_8_n_307) & (mul_22_8_n_370 | mul_22_8_n_103));
 assign mul_22_8_n_543 = ~((mul_22_8_n_237 | mul_22_8_n_75) & (mul_22_8_n_371 | mul_22_8_n_186));
 assign mul_22_8_n_542 = ~((mul_22_8_n_232 | mul_22_8_n_73) & (mul_22_8_n_366 | mul_22_8_n_187));
 assign mul_22_8_n_541 = ~((mul_22_8_n_233 | mul_22_8_n_179) & (mul_22_8_n_367 | mul_22_8_n_161));
 assign mul_22_8_n_540 = ~((mul_22_8_n_232 | mul_22_8_n_265) & (mul_22_8_n_366 | mul_22_8_n_264));
 assign mul_22_8_n_539 = ~((mul_22_8_n_235 | mul_22_8_n_144) & (mul_22_8_n_369 | mul_22_8_n_130));
 assign mul_22_8_n_538 = ~((mul_22_8_n_237 | mul_22_8_n_281) & (mul_22_8_n_371 | mul_22_8_n_282));
 assign mul_22_8_n_537 = ~((mul_22_8_n_236 | mul_22_8_n_267) & (mul_22_8_n_370 | mul_22_8_n_292));
 assign mul_22_8_n_536 = ~((mul_22_8_n_234 | mul_22_8_n_99) & (mul_22_8_n_368 | mul_22_8_n_96));
 assign mul_22_8_n_535 = ~((mul_22_8_n_240 | mul_22_8_n_156) & (mul_22_8_n_374 | mul_22_8_n_157));
 assign mul_22_8_n_534 = ~((mul_22_8_n_235 | mul_22_8_n_163) & (mul_22_8_n_369 | mul_22_8_n_164));
 assign mul_22_8_n_533 = ~((mul_22_8_n_238 | mul_22_8_n_145) & (mul_22_8_n_372 | mul_22_8_n_146));
 assign mul_22_8_n_532 = ~((mul_22_8_n_234 | mul_22_8_n_291) & (mul_22_8_n_368 | mul_22_8_n_290));
 assign mul_22_8_n_531 = ~((mul_22_8_n_235 | mul_22_8_n_183) & (mul_22_8_n_369 | mul_22_8_n_184));
 assign mul_22_8_n_530 = ~((mul_22_8_n_238 | mul_22_8_n_169) & (mul_22_8_n_372 | mul_22_8_n_170));
 assign mul_22_8_n_529 = ~((mul_22_8_n_239 | mul_22_8_n_132) & (mul_22_8_n_373 | mul_22_8_n_131));
 assign mul_22_8_n_528 = ~((mul_22_8_n_236 | mul_22_8_n_149) & (mul_22_8_n_370 | mul_22_8_n_191));
 assign mul_22_8_n_527 = ~((mul_22_8_n_235 | mul_22_8_n_184) & (mul_22_8_n_369 | mul_22_8_n_163));
 assign mul_22_8_n_526 = ~((mul_22_8_n_233 | mul_22_8_n_301) & (mul_22_8_n_367 | mul_22_8_n_357));
 assign mul_22_8_n_525 = ~((mul_22_8_n_240 | mul_22_8_n_105) & (mul_22_8_n_374 | mul_22_8_n_104));
 assign mul_22_8_n_524 = ~((mul_22_8_n_241 | mul_22_8_n_79) & (mul_22_8_n_375 | mul_22_8_n_80));
 assign mul_22_8_n_523 = ~((mul_22_8_n_237 | mul_22_8_n_125) & (mul_22_8_n_371 | mul_22_8_n_124));
 assign mul_22_8_n_522 = ~((mul_22_8_n_233 | mul_22_8_n_311) & (mul_22_8_n_367 | mul_22_8_n_312));
 assign mul_22_8_n_521 = ~((mul_22_8_n_236 | mul_22_8_n_292) & (mul_22_8_n_370 | mul_22_8_n_307));
 assign mul_22_8_n_520 = ~((mul_22_8_n_238 | mul_22_8_n_146) & (mul_22_8_n_372 | mul_22_8_n_127));
 assign mul_22_8_n_519 = ~((mul_22_8_n_232 | mul_22_8_n_168) & (mul_22_8_n_366 | mul_22_8_n_167));
 assign mul_22_8_n_518 = ~((mul_22_8_n_233 | mul_22_8_n_336) & (mul_22_8_n_367 | mul_22_8_n_137));
 assign mul_22_8_n_517 = ~((mul_22_8_n_238 | mul_22_8_n_153) & (mul_22_8_n_372 | mul_22_8_n_200));
 assign mul_22_8_n_516 = ~((mul_22_8_n_233 | mul_22_8_n_333) & (mul_22_8_n_367 | mul_22_8_n_336));
 assign mul_22_8_n_515 = ~((mul_22_8_n_233 | mul_22_8_n_261) & (mul_22_8_n_367 | mul_22_8_n_333));
 assign mul_22_8_n_514 = ~((mul_22_8_n_241 | mul_22_8_n_89) & (mul_22_8_n_375 | mul_22_8_n_88));
 assign mul_22_8_n_513 = ~((mul_22_8_n_232 | mul_22_8_n_188) & (mul_22_8_n_366 | mul_22_8_n_168));
 assign mul_22_8_n_512 = ~((mul_22_8_n_235 | mul_22_8_n_322) & (mul_22_8_n_369 | mul_22_8_n_306));
 assign mul_22_8_n_511 = ~((mul_22_8_n_241 | mul_22_8_n_138) & (mul_22_8_n_375 | mul_22_8_n_114));
 assign mul_22_8_n_510 = ~((mul_22_8_n_233 | mul_22_8_n_180) & (mul_22_8_n_367 | mul_22_8_n_179));
 assign mul_22_8_n_509 = ~((mul_22_8_n_240 | mul_22_8_n_93) & (mul_22_8_n_374 | mul_22_8_n_94));
 assign mul_22_8_n_508 = ~((mul_22_8_n_232 | mul_22_8_n_332) & (mul_22_8_n_366 | mul_22_8_n_330));
 assign mul_22_8_n_507 = ~((mul_22_8_n_234 | mul_22_8_n_310) & (mul_22_8_n_368 | mul_22_8_n_291));
 assign mul_22_8_n_506 = ~((mul_22_8_n_241 | mul_22_8_n_102) & (mul_22_8_n_375 | mul_22_8_n_101));
 assign mul_22_8_n_505 = ~((mul_22_8_n_237 | mul_22_8_n_258) & (mul_22_8_n_371 | mul_22_8_n_259));
 assign mul_22_8_n_504 = ~((mul_22_8_n_240 | mul_22_8_n_120) & (mul_22_8_n_374 | mul_22_8_n_105));
 assign mul_22_8_n_503 = ~((mul_22_8_n_234 | mul_22_8_n_346) & (mul_22_8_n_368 | mul_22_8_n_99));
 assign mul_22_8_n_502 = ~((mul_22_8_n_241 | mul_22_8_n_88) & (mul_22_8_n_375 | mul_22_8_n_79));
 assign mul_22_8_n_501 = ~((mul_22_8_n_235 | mul_22_8_n_204) & (mul_22_8_n_369 | mul_22_8_n_183));
 assign mul_22_8_n_500 = ~((mul_22_8_n_237 | mul_22_8_n_74) & (mul_22_8_n_371 | mul_22_8_n_75));
 assign mul_22_8_n_499 = ~((mul_22_8_n_233 | mul_22_8_n_327) & (mul_22_8_n_367 | mul_22_8_n_311));
 assign mul_22_8_n_498 = ~((mul_22_8_n_242 | mul_22_8_n_90) & (mul_22_8_n_376 | mul_22_8_n_100));
 assign mul_22_8_n_497 = ~((mul_22_8_n_237 | mul_22_8_n_342) & (mul_22_8_n_371 | mul_22_8_n_74));
 assign mul_22_8_n_496 = ~((mul_22_8_n_236 | mul_22_8_n_173) & (mul_22_8_n_370 | mul_22_8_n_149));
 assign mul_22_8_n_495 = ~((mul_22_8_n_237 | mul_22_8_n_141) & (mul_22_8_n_371 | mul_22_8_n_125));
 assign mul_22_8_n_494 = ~((mul_22_8_n_233 | mul_22_8_n_202) & (mul_22_8_n_367 | mul_22_8_n_203));
 assign mul_22_8_n_493 = ~((mul_22_8_n_0 | mul_22_8_n_166) & (mul_22_8_n_378 | mul_22_8_n_177));
 assign mul_22_8_n_492 = ~((mul_22_8_n_232 | mul_22_8_n_189) & (mul_22_8_n_366 | mul_22_8_n_70));
 assign mul_22_8_n_491 = ~((mul_22_8_n_239 | mul_22_8_n_118) & (mul_22_8_n_373 | mul_22_8_n_117));
 assign mul_22_8_n_490 = ~((mul_22_8_n_234 | mul_22_8_n_171) & (mul_22_8_n_368 | mul_22_8_n_155));
 assign mul_22_8_n_489 = ~((mul_22_8_n_239 | mul_22_8_n_76) & (mul_22_8_n_373 | mul_22_8_n_78));
 assign mul_22_8_n_488 = ~((mul_22_8_n_234 | mul_22_8_n_309) & (mul_22_8_n_368 | mul_22_8_n_310));
 assign mul_22_8_n_487 = ~((mul_22_8_n_238 | mul_22_8_n_200) & (mul_22_8_n_372 | mul_22_8_n_201));
 assign mul_22_8_n_486 = ~((mul_22_8_n_242 | mul_22_8_n_84) & (mul_22_8_n_376 | mul_22_8_n_83));
 assign mul_22_8_n_485 = ~((mul_22_8_n_235 | mul_22_8_n_288) & (mul_22_8_n_369 | mul_22_8_n_289));
 assign mul_22_8_n_484 = ~((mul_22_8_n_240 | mul_22_8_n_119) & (mul_22_8_n_374 | mul_22_8_n_120));
 assign mul_22_8_n_483 = ~((mul_22_8_n_234 | mul_22_8_n_344) & (mul_22_8_n_368 | mul_22_8_n_346));
 assign mul_22_8_n_482 = ~((mul_22_8_n_236 | mul_22_8_n_266) & (mul_22_8_n_370 | mul_22_8_n_267));
 assign mul_22_8_n_481 = ~((mul_22_8_n_238 | mul_22_8_n_115) & (mul_22_8_n_372 | mul_22_8_n_116));
 assign mul_22_8_n_480 = ~((mul_22_8_n_242 | mul_22_8_n_91) & (mul_22_8_n_376 | mul_22_8_n_90));
 assign mul_22_8_n_479 = ~((mul_22_8_n_233 | mul_22_8_n_328) & (mul_22_8_n_367 | mul_22_8_n_327));
 assign mul_22_8_n_478 = ~((mul_22_8_n_237 | mul_22_8_n_339) & (mul_22_8_n_371 | mul_22_8_n_342));
 assign mul_22_8_n_477 = ~((mul_22_8_n_232 | mul_22_8_n_167) & (mul_22_8_n_366 | mul_22_8_n_152));
 assign mul_22_8_n_476 = ~((mul_22_8_n_232 | mul_22_8_n_280) & (mul_22_8_n_366 | mul_22_8_n_279));
 assign mul_22_8_n_475 = ~((mul_22_8_n_234 | mul_22_8_n_326) & (mul_22_8_n_368 | mul_22_8_n_309));
 assign mul_22_8_n_474 = ~((mul_22_8_n_235 | mul_22_8_n_205) & (mul_22_8_n_369 | mul_22_8_n_204));
 assign mul_22_8_n_473 = ~((mul_22_8_n_239 | mul_22_8_n_150) & (mul_22_8_n_373 | mul_22_8_n_151));
 assign mul_22_8_n_472 = ~((mul_22_8_n_236 | mul_22_8_n_174) & (mul_22_8_n_370 | mul_22_8_n_173));
 assign mul_22_8_n_471 = ~((mul_22_8_n_234 | mul_22_8_n_257) & (mul_22_8_n_368 | mul_22_8_n_256));
 assign mul_22_8_n_470 = ~((mul_22_8_n_237 | mul_22_8_n_142) & (mul_22_8_n_371 | mul_22_8_n_141));
 assign mul_22_8_n_469 = ~((mul_22_8_n_234 | mul_22_8_n_273) & (mul_22_8_n_368 | mul_22_8_n_274));
 assign mul_22_8_n_468 = ~((mul_22_8_n_233 | mul_22_8_n_294) & (mul_22_8_n_367 | mul_22_8_n_293));
 assign mul_22_8_n_467 = ~((mul_22_8_n_232 | mul_22_8_n_308) & (mul_22_8_n_366 | mul_22_8_n_341));
 assign mul_22_8_n_466 = ~((mul_22_8_n_234 | mul_22_8_n_274) & (mul_22_8_n_368 | mul_22_8_n_257));
 assign mul_22_8_n_465 = ~((mul_22_8_n_239 | mul_22_8_n_182) & (mul_22_8_n_373 | mul_22_8_n_181));
 assign mul_22_8_n_464 = ~((mul_22_8_n_239 | mul_22_8_n_181) & (mul_22_8_n_373 | mul_22_8_n_150));
 assign mul_22_8_n_463 = ~((mul_22_8_n_235 | mul_22_8_n_305) & (mul_22_8_n_369 | mul_22_8_n_288));
 assign mul_22_8_n_462 = ~((mul_22_8_n_234 | mul_22_8_n_172) & (mul_22_8_n_368 | mul_22_8_n_171));
 assign mul_22_8_n_461 = ~((mul_22_8_n_240 | mul_22_8_n_134) & (mul_22_8_n_374 | mul_22_8_n_119));
 assign mul_22_8_n_460 = ~((mul_22_8_n_241 | mul_22_8_n_101) & (mul_22_8_n_375 | mul_22_8_n_89));
 assign mul_22_8_n_459 = ~((mul_22_8_n_235 | mul_22_8_n_148) & (mul_22_8_n_369 | mul_22_8_n_205));
 assign mul_22_8_n_458 = ~((mul_22_8_n_235 | mul_22_8_n_143) & (mul_22_8_n_369 | mul_22_8_n_144));
 assign mul_22_8_n_457 = ~((mul_22_8_n_236 | mul_22_8_n_287) & (mul_22_8_n_370 | mul_22_8_n_266));
 assign mul_22_8_n_456 = ~((mul_22_8_n_242 | mul_22_8_n_82) & (mul_22_8_n_376 | mul_22_8_n_91));
 assign mul_22_8_n_455 = ~((mul_22_8_n_233 | mul_22_8_n_270) & (mul_22_8_n_367 | mul_22_8_n_328));
 assign mul_22_8_n_454 = ~((mul_22_8_n_237 | mul_22_8_n_185) & (mul_22_8_n_371 | mul_22_8_n_160));
 assign mul_22_8_n_453 = ~((mul_22_8_n_233 | mul_22_8_n_260) & (mul_22_8_n_367 | mul_22_8_n_261));
 assign mul_22_8_n_452 = ~((mul_22_8_n_238 | mul_22_8_n_252) & (mul_22_8_n_372 | mul_22_8_n_253));
 assign mul_22_8_n_451 = ~((mul_22_8_n_239 | mul_22_8_n_107) & (mul_22_8_n_373 | mul_22_8_n_95));
 assign mul_22_8_n_450 = ~((mul_22_8_n_232 | mul_22_8_n_295) & (mul_22_8_n_366 | mul_22_8_n_280));
 assign mul_22_8_n_449 = ~((mul_22_8_n_233 | mul_22_8_n_293) & (mul_22_8_n_367 | mul_22_8_n_278));
 assign mul_22_8_n_448 = ~((mul_22_8_n_234 | mul_22_8_n_325) & (mul_22_8_n_368 | mul_22_8_n_326));
 assign mul_22_8_n_447 = ~((mul_22_8_n_238 | mul_22_8_n_140) & (mul_22_8_n_372 | mul_22_8_n_153));
 assign mul_22_8_n_446 = ~((mul_22_8_n_238 | mul_22_8_n_116) & (mul_22_8_n_372 | mul_22_8_n_108));
 assign mul_22_8_n_445 = ~((mul_22_8_n_233 | mul_22_8_n_277) & (mul_22_8_n_367 | mul_22_8_n_260));
 assign mul_22_8_n_444 = ~((mul_22_8_n_235 | mul_22_8_n_306) & (mul_22_8_n_369 | mul_22_8_n_305));
 assign mul_22_8_n_443 = ~((mul_22_8_n_240 | mul_22_8_n_190) & (mul_22_8_n_374 | mul_22_8_n_156));
 assign mul_22_8_n_442 = ~((mul_22_8_n_240 | mul_22_8_n_133) & (mul_22_8_n_374 | mul_22_8_n_134));
 assign mul_22_8_n_441 = ~((mul_22_8_n_236 | mul_22_8_n_198) & (mul_22_8_n_370 | mul_22_8_n_174));
 assign mul_22_8_n_562 = ~((mul_22_8_n_363 & mul_22_8_n_340) | (mul_22_8_n_365 & mul_22_8_n_331));
 assign mul_22_8_n_561 = ((mul_22_8_n_232 | mul_22_8_n_165) & (mul_22_8_n_366 | mul_22_8_n_189));
 assign mul_22_8_n_560 = ((mul_22_8_n_232 | mul_22_8_n_302) & (mul_22_8_n_366 | mul_22_8_n_308));
 assign mul_22_8_n_559 = ~((mul_22_8_n_363 & mul_22_8_n_71) | (mul_22_8_n_365 & mul_22_8_n_72));
 assign mul_22_8_n_558 = ~((mul_22_8_n_232 | mul_22_8_n_330) & (mul_22_8_n_366 | mul_22_8_n_329));
 assign mul_22_8_n_437 = ~((mul_22_8_n_316 | mul_22_8_n_34) & (mul_22_8_n_362 | mul_22_8_n_297));
 assign mul_22_8_n_436 = ~(({in2[12]} & {in1[0]}) | ({in2[11]} & ({in2[12]} ^ {in1[0]})));
 assign mul_22_8_n_435 = ~(({in2[4]} & {in1[0]}) | ({in2[3]} & ({in2[4]} ^ {in1[0]})));
 assign mul_22_8_n_434 = ~(({in2[24]} & {in1[0]}) | ({in2[23]} & ({in2[24]} ^ {in1[0]})));
 assign mul_22_8_n_433 = ~(({in2[20]} & {in1[0]}) | ({in2[19]} & ({in2[20]} ^ {in1[0]})));
 assign mul_22_8_n_432 = ~(({in2[8]} & {in1[0]}) | ({in2[7]} & ({in2[8]} ^ {in1[0]})));
 assign mul_22_8_n_431 = ~(({in2[14]} & {in1[0]}) | ({in2[13]} & ({in2[14]} ^ {in1[0]})));
 assign mul_22_8_n_430 = ~(({in2[30]} & {in1[0]}) | ({in2[29]} & ({in2[30]} ^ {in1[0]})));
 assign mul_22_8_n_429 = ~(({in2[28]} & {in1[0]}) | ({in2[27]} & ({in2[28]} ^ {in1[0]})));
 assign mul_22_8_n_428 = ~(({in2[22]} & {in1[0]}) | ({in2[21]} & ({in2[22]} ^ {in1[0]})));
 assign mul_22_8_n_427 = ~(({in2[2]} & {in1[0]}) | ({in2[1]} & ({in2[2]} ^ {in1[0]})));
 assign mul_22_8_n_426 = ~(({in2[26]} & {in1[0]}) | ({in2[25]} & ({in2[26]} ^ {in1[0]})));
 assign mul_22_8_n_425 = ~(({in2[6]} & {in1[0]}) | ({in2[5]} & ({in2[6]} ^ {in1[0]})));
 assign mul_22_8_n_424 = ~(({in2[10]} & {in1[0]}) | ({in2[9]} & ({in2[10]} ^ {in1[0]})));
 assign mul_22_8_n_423 = ~(({in2[16]} & {in1[0]}) | ({in2[15]} & ({in2[16]} ^ {in1[0]})));
 assign mul_22_8_n_422 = ~(({in2[18]} & {in1[0]}) | ({in2[17]} & ({in2[18]} ^ {in1[0]})));
 assign mul_22_8_n_421 = ~((mul_22_8_n_196 | mul_22_8_n_34) & (mul_22_8_n_362 | mul_22_8_n_175));
 assign mul_22_8_n_420 = ~((mul_22_8_n_352 | mul_22_8_n_34) & (mul_22_8_n_362 | mul_22_8_n_338));
 assign mul_22_8_n_419 = ~((mul_22_8_n_347 | mul_22_8_n_34) & (mul_22_8_n_362 | mul_22_8_n_358));
 assign mul_22_8_n_440 = ~((mul_22_8_n_158 & {in2[0]}) | (mul_22_8_n_361 & mul_22_8_n_55));
 assign mul_22_8_n_418 = ~((mul_22_8_n_218 & {in2[0]}) | (mul_22_8_n_361 & mul_22_8_n_353));
 assign mul_22_8_n_439 = ~((mul_22_8_n_197 & {in2[0]}) | (mul_22_8_n_361 & mul_22_8_n_195));
 assign mul_22_8_n_438 = ~((mul_22_8_n_268 & {in2[0]}) | (mul_22_8_n_361 & mul_22_8_n_269));
 assign mul_22_8_n_410 = ~((mul_22_8_n_356 | mul_22_8_n_34) & (mul_22_8_n_362 | mul_22_8_n_351));
 assign mul_22_8_n_409 = ~((mul_22_8_n_334 | mul_22_8_n_34) & (mul_22_8_n_362 | mul_22_8_n_315));
 assign mul_22_8_n_408 = ~((mul_22_8_n_349 | mul_22_8_n_34) & (mul_22_8_n_362 | mul_22_8_n_317));
 assign mul_22_8_n_407 = ~((mul_22_8_n_345 | mul_22_8_n_34) & (mul_22_8_n_362 | mul_22_8_n_255));
 assign mul_22_8_n_406 = ~((mul_22_8_n_255 | mul_22_8_n_34) & (mul_22_8_n_362 | mul_22_8_n_349));
 assign mul_22_8_n_405 = ((mul_22_8_n_269 & {in2[0]}) | (mul_22_8_n_361 & mul_22_8_n_247));
 assign mul_22_8_n_404 = ~((mul_22_8_n_335 | mul_22_8_n_34) & (mul_22_8_n_362 | mul_22_8_n_334));
 assign mul_22_8_n_403 = ~((mul_22_8_n_299 | mul_22_8_n_34) & (mul_22_8_n_362 | mul_22_8_n_285));
 assign mul_22_8_n_402 = ~((mul_22_8_n_249 | mul_22_8_n_34) & (mul_22_8_n_362 | mul_22_8_n_356));
 assign mul_22_8_n_401 = ~((mul_22_8_n_248 | mul_22_8_n_34) & (mul_22_8_n_362 | mul_22_8_n_249));
 assign mul_22_8_n_400 = ~((mul_22_8_n_351 | mul_22_8_n_34) & (mul_22_8_n_362 | mul_22_8_n_86));
 assign mul_22_8_n_399 = ~((mul_22_8_n_358 | mul_22_8_n_34) & (mul_22_8_n_362 | mul_22_8_n_345));
 assign mul_22_8_n_398 = ~((mul_22_8_n_337 | mul_22_8_n_34) & (mul_22_8_n_362 | mul_22_8_n_335));
 assign mul_22_8_n_397 = ((mul_22_8_n_92 & {in2[0]}) | (mul_22_8_n_361 & mul_22_8_n_197));
 assign mul_22_8_n_396 = ((mul_22_8_n_283 & {in2[0]}) | (mul_22_8_n_361 & mul_22_8_n_268));
 assign mul_22_8_n_395 = ~((mul_22_8_n_317 | mul_22_8_n_34) & (mul_22_8_n_362 | mul_22_8_n_337));
 assign mul_22_8_n_417 = ~((mul_22_8_n_176 & {in2[0]}) | (mul_22_8_n_361 & mul_22_8_n_158));
 assign mul_22_8_n_416 = ~((mul_22_8_n_284 & {in2[0]}) | (mul_22_8_n_361 & mul_22_8_n_283));
 assign mul_22_8_n_415 = ((mul_22_8_n_315 | mul_22_8_n_34) & (mul_22_8_n_362 | mul_22_8_n_316));
 assign mul_22_8_n_414 = ~((~mul_22_8_n_297 & ~mul_22_8_n_34) | (mul_22_8_n_361 & mul_22_8_n_298));
 assign mul_22_8_n_413 = ~((~mul_22_8_n_175 & ~mul_22_8_n_34) | (mul_22_8_n_361 & mul_22_8_n_176));
 assign mul_22_8_n_412 = ~((mul_22_8_n_87 & {in2[0]}) | (mul_22_8_n_361 & mul_22_8_n_92));
 assign mul_22_8_n_411 = ((mul_22_8_n_338 | mul_22_8_n_34) & (mul_22_8_n_362 | mul_22_8_n_347));
 assign mul_22_8_n_393 = ~(n_155 | mul_22_8_n_9);
 assign mul_22_8_n_392 = ~(mul_22_8_n_244 | mul_22_8_n_9);
 assign mul_22_8_n_391 = ~(mul_22_8_n_233 | mul_22_8_n_9);
 assign mul_22_8_n_390 = ~(mul_22_8_n_240 | mul_22_8_n_9);
 assign mul_22_8_n_389 = ~(mul_22_8_n_241 | mul_22_8_n_9);
 assign mul_22_8_n_388 = ~(mul_22_8_n_236 | mul_22_8_n_9);
 assign mul_22_8_n_387 = ~(mul_22_8_n_238 | mul_22_8_n_9);
 assign mul_22_8_n_386 = ~(mul_22_8_n_237 | mul_22_8_n_9);
 assign mul_22_8_n_385 = ~(mul_22_8_n_234 | mul_22_8_n_9);
 assign mul_22_8_n_384 = ~(mul_22_8_n_235 | mul_22_8_n_9);
 assign mul_22_8_n_383 = ~(mul_22_8_n_242 | mul_22_8_n_9);
 assign mul_22_8_n_382 = (mul_22_8_n_245 & {in1[0]});
 assign mul_22_8_n_381 = ~(mul_22_8_n_239 | mul_22_8_n_9);
 assign mul_22_8_n_380 = ~(mul_22_8_n_0 | mul_22_8_n_9);
 assign mul_22_8_n_394 = ~(mul_22_8_n_363 & {in1[0]});
 assign mul_22_8_n_365 = ~mul_22_8_n_366;
 assign mul_22_8_n_364 = ~(mul_22_8_n_245 & (mul_22_8_n_48 | (mul_22_8_n_35 & {in2[31]})));
 assign mul_22_8_n_379 = ~(mul_22_8_n_244 & (mul_22_8_n_49 | (mul_22_8_n_25 & {in2[28]})));
 assign mul_22_8_n_378 = ~(mul_22_8_n_0 & (mul_22_8_n_50 | (mul_22_8_n_21 & {in2[26]})));
 assign mul_22_8_n_377 = ~(n_155 & mul_22_8_n_211);
 assign mul_22_8_n_376 = ~(mul_22_8_n_242 & mul_22_8_n_212);
 assign mul_22_8_n_375 = ~(mul_22_8_n_241 & mul_22_8_n_215);
 assign mul_22_8_n_374 = ~(mul_22_8_n_240 & mul_22_8_n_216);
 assign mul_22_8_n_373 = ~(mul_22_8_n_239 & mul_22_8_n_217);
 assign mul_22_8_n_372 = ~(mul_22_8_n_238 & mul_22_8_n_231);
 assign mul_22_8_n_371 = ~(mul_22_8_n_237 & mul_22_8_n_219);
 assign mul_22_8_n_370 = ~(mul_22_8_n_236 & mul_22_8_n_220);
 assign mul_22_8_n_369 = ~(mul_22_8_n_235 & mul_22_8_n_221);
 assign mul_22_8_n_368 = ~(mul_22_8_n_234 & mul_22_8_n_224);
 assign mul_22_8_n_367 = ~(mul_22_8_n_233 & mul_22_8_n_227);
 assign mul_22_8_n_366 = ~(mul_22_8_n_232 & mul_22_8_n_228);
 assign mul_22_8_n_363 = ~mul_22_8_n_232;
 assign mul_22_8_n_361 = ~mul_22_8_n_362;
 assign mul_22_8_n_362 = ~({in2[1]} & mul_22_8_n_34);
 assign mul_22_8_n_353 = ~mul_22_8_n_352;
 assign mul_22_8_n_341 = ~mul_22_8_n_340;
 assign mul_22_8_n_332 = ~mul_22_8_n_331;
 assign mul_22_8_n_299 = ~mul_22_8_n_298;
 assign mul_22_8_n_285 = ~mul_22_8_n_284;
 assign mul_22_8_n_248 = ~mul_22_8_n_247;
 assign mul_22_8_n_231 = ~((mul_22_8_n_11 & ~{in2[14]}) | ({in2[15]} & {in2[14]}));
 assign mul_22_8_n_230 = ~((mul_22_8_n_9 & {in2[25]}) | (mul_22_8_n_18 & {in1[0]}));
 assign mul_22_8_n_229 = ~(({in2[3]} & ~{in1[29]}) | (mul_22_8_n_29 & {in1[29]}));
 assign mul_22_8_n_228 = ~((mul_22_8_n_29 & ~{in2[2]}) | ({in2[3]} & {in2[2]}));
 assign mul_22_8_n_227 = ~((mul_22_8_n_30 & ~{in2[4]}) | ({in2[5]} & {in2[4]}));
 assign mul_22_8_n_226 = ~(({in1[0]} & ~{in2[31]}) | (mul_22_8_n_9 & {in2[31]}));
 assign mul_22_8_n_225 = ~(({in2[5]} & ~{in1[27]}) | (mul_22_8_n_30 & {in1[27]}));
 assign mul_22_8_n_224 = ~((mul_22_8_n_31 & ~{in2[6]}) | ({in2[7]} & {in2[6]}));
 assign mul_22_8_n_223 = ~(({in2[7]} & ~{in1[25]}) | (mul_22_8_n_31 & {in1[25]}));
 assign mul_22_8_n_222 = ~(({in2[9]} & ~{in1[23]}) | (mul_22_8_n_32 & {in1[23]}));
 assign mul_22_8_n_221 = ~((mul_22_8_n_32 & ~{in2[8]}) | ({in2[9]} & {in2[8]}));
 assign mul_22_8_n_220 = ~((mul_22_8_n_33 & ~{in2[10]}) | ({in2[11]} & {in2[10]}));
 assign mul_22_8_n_219 = ~((mul_22_8_n_10 & ~{in2[12]}) | ({in2[13]} & {in2[12]}));
 assign mul_22_8_n_218 = ~((mul_22_8_n_8 & ~{in1[31]}) | ({in2[1]} & {in1[31]}));
 assign mul_22_8_n_217 = ~((mul_22_8_n_12 & ~{in2[16]}) | ({in2[17]} & {in2[16]}));
 assign mul_22_8_n_216 = ~((mul_22_8_n_13 & ~{in2[18]}) | ({in2[19]} & {in2[18]}));
 assign mul_22_8_n_215 = ~((mul_22_8_n_36 & ~{in2[20]}) | ({in2[21]} & {in2[20]}));
 assign mul_22_8_n_214 = ~((mul_22_8_n_27 & {in2[11]}) | (mul_22_8_n_33 & {in1[21]}));
 assign mul_22_8_n_213 = ~((mul_22_8_n_44 & {in2[17]}) | (mul_22_8_n_12 & {in1[15]}));
 assign mul_22_8_n_212 = ~((mul_22_8_n_17 & ~{in2[22]}) | ({in2[23]} & {in2[22]}));
 assign mul_22_8_n_211 = ~((mul_22_8_n_18 & ~{in2[24]}) | ({in2[25]} & {in2[24]}));
 assign mul_22_8_n_210 = ~((mul_22_8_n_9 & {in2[29]}) | (mul_22_8_n_25 & {in1[0]}));
 assign mul_22_8_n_209 = ~((mul_22_8_n_45 & {in2[13]}) | (mul_22_8_n_10 & {in1[19]}));
 assign mul_22_8_n_208 = ~((mul_22_8_n_23 & {in2[15]}) | (mul_22_8_n_11 & {in1[17]}));
 assign mul_22_8_n_207 = ~((mul_22_8_n_9 & {in2[27]}) | (mul_22_8_n_21 & {in1[0]}));
 assign mul_22_8_n_206 = ~((mul_22_8_n_14 & {in2[29]}) | (mul_22_8_n_25 & {in1[3]}));
 assign mul_22_8_n_360 = ~({in2[1]} & ~asc001_0_);
 assign mul_22_8_n_359 = ~(({in2[5]} & ~{in1[23]}) | (mul_22_8_n_30 & {in1[23]}));
 assign mul_22_8_n_358 = ~(({in2[1]} & ~{in1[27]}) | (mul_22_8_n_8 & {in1[27]}));
 assign mul_22_8_n_357 = ~(({in2[5]} & ~{in1[25]}) | (mul_22_8_n_30 & {in1[25]}));
 assign mul_22_8_n_356 = ~((mul_22_8_n_40 & {in2[1]}) | (mul_22_8_n_8 & {in1[9]}));
 assign mul_22_8_n_355 = ~(({in2[7]} & ~{in1[22]}) | (mul_22_8_n_31 & {in1[22]}));
 assign mul_22_8_n_354 = ~(({in2[7]} & ~{in1[23]}) | (mul_22_8_n_31 & {in1[23]}));
 assign mul_22_8_n_352 = ~(({in2[1]} & ~{in1[30]}) | (mul_22_8_n_8 & {in1[30]}));
 assign mul_22_8_n_351 = ~((mul_22_8_n_41 & {in2[1]}) | (mul_22_8_n_8 & {in1[8]}));
 assign mul_22_8_n_350 = ~(({in2[7]} & ~{in1[24]}) | (mul_22_8_n_31 & {in1[24]}));
 assign mul_22_8_n_349 = ~(({in2[1]} & ~{in1[24]}) | (mul_22_8_n_8 & {in1[24]}));
 assign mul_22_8_n_348 = ~(({in2[9]} & ~{in1[22]}) | (mul_22_8_n_32 & {in1[22]}));
 assign mul_22_8_n_347 = ~(({in2[1]} & ~{in1[28]}) | (mul_22_8_n_8 & {in1[28]}));
 assign mul_22_8_n_346 = ~((mul_22_8_n_19 & {in2[7]}) | (mul_22_8_n_31 & {in1[10]}));
 assign mul_22_8_n_345 = ~(({in2[1]} & ~{in1[26]}) | (mul_22_8_n_8 & {in1[26]}));
 assign mul_22_8_n_344 = ~((mul_22_8_n_42 & {in2[7]}) | (mul_22_8_n_31 & {in1[11]}));
 assign mul_22_8_n_343 = ~((mul_22_8_n_42 & {in2[9]}) | (mul_22_8_n_32 & {in1[11]}));
 assign mul_22_8_n_342 = ~((mul_22_8_n_43 & {in2[13]}) | (mul_22_8_n_10 & {in1[12]}));
 assign mul_22_8_n_340 = ~((mul_22_8_n_29 & ~{in1[23]}) | ({in2[3]} & {in1[23]}));
 assign mul_22_8_n_339 = ~((mul_22_8_n_20 & {in2[13]}) | (mul_22_8_n_10 & {in1[13]}));
 assign mul_22_8_n_338 = ~(({in2[1]} & ~{in1[29]}) | (mul_22_8_n_8 & {in1[29]}));
 assign mul_22_8_n_337 = ~(({in2[1]} & ~{in1[22]}) | (mul_22_8_n_8 & {in1[22]}));
 assign mul_22_8_n_336 = ~((mul_22_8_n_19 & {in2[5]}) | (mul_22_8_n_30 & {in1[10]}));
 assign mul_22_8_n_335 = ~((mul_22_8_n_27 & {in2[1]}) | (mul_22_8_n_8 & {in1[21]}));
 assign mul_22_8_n_334 = ~((mul_22_8_n_46 & {in2[1]}) | (mul_22_8_n_8 & {in1[20]}));
 assign mul_22_8_n_333 = ~((mul_22_8_n_42 & {in2[5]}) | (mul_22_8_n_30 & {in1[11]}));
 assign mul_22_8_n_331 = ~((mul_22_8_n_29 & ~{in1[22]}) | ({in2[3]} & {in1[22]}));
 assign mul_22_8_n_330 = ~((mul_22_8_n_27 & {in2[3]}) | (mul_22_8_n_29 & {in1[21]}));
 assign mul_22_8_n_329 = ~((mul_22_8_n_46 & {in2[3]}) | (mul_22_8_n_29 & {in1[20]}));
 assign mul_22_8_n_328 = ~((mul_22_8_n_27 & {in2[5]}) | (mul_22_8_n_30 & {in1[21]}));
 assign mul_22_8_n_327 = ~((mul_22_8_n_46 & {in2[5]}) | (mul_22_8_n_30 & {in1[20]}));
 assign mul_22_8_n_326 = ~((mul_22_8_n_46 & {in2[7]}) | (mul_22_8_n_31 & {in1[20]}));
 assign mul_22_8_n_325 = ~((mul_22_8_n_27 & {in2[7]}) | (mul_22_8_n_31 & {in1[21]}));
 assign mul_22_8_n_324 = ~((mul_22_8_n_22 & {in2[17]}) | (mul_22_8_n_12 & {in1[14]}));
 assign mul_22_8_n_323 = ~(({in2[3]} & ~{in1[27]}) | (mul_22_8_n_29 & {in1[27]}));
 assign mul_22_8_n_322 = ~((mul_22_8_n_46 & {in2[9]}) | (mul_22_8_n_32 & {in1[20]}));
 assign mul_22_8_n_321 = ~((mul_22_8_n_27 & {in2[9]}) | (mul_22_8_n_32 & {in1[21]}));
 assign mul_22_8_n_320 = ~(({in2[3]} & ~{in1[26]}) | (mul_22_8_n_29 & {in1[26]}));
 assign mul_22_8_n_319 = ~((mul_22_8_n_46 & {in2[11]}) | (mul_22_8_n_33 & {in1[20]}));
 assign mul_22_8_n_318 = ~(({in2[3]} & ~{in1[28]}) | (mul_22_8_n_29 & {in1[28]}));
 assign mul_22_8_n_317 = ~(({in2[1]} & ~{in1[23]}) | (mul_22_8_n_8 & {in1[23]}));
 assign mul_22_8_n_316 = ~((mul_22_8_n_26 & {in2[1]}) | (mul_22_8_n_8 & {in1[18]}));
 assign mul_22_8_n_315 = ~((mul_22_8_n_45 & {in2[1]}) | (mul_22_8_n_8 & {in1[19]}));
 assign mul_22_8_n_314 = ~((mul_22_8_n_45 & {in2[3]}) | (mul_22_8_n_29 & {in1[19]}));
 assign mul_22_8_n_313 = ~((mul_22_8_n_26 & {in2[3]}) | (mul_22_8_n_29 & {in1[18]}));
 assign mul_22_8_n_312 = ~((mul_22_8_n_26 & {in2[5]}) | (mul_22_8_n_30 & {in1[18]}));
 assign mul_22_8_n_311 = ~((mul_22_8_n_45 & {in2[5]}) | (mul_22_8_n_30 & {in1[19]}));
 assign mul_22_8_n_310 = ~((mul_22_8_n_26 & {in2[7]}) | (mul_22_8_n_31 & {in1[18]}));
 assign mul_22_8_n_309 = ~((mul_22_8_n_45 & {in2[7]}) | (mul_22_8_n_31 & {in1[19]}));
 assign mul_22_8_n_308 = ~(({in2[3]} & ~{in1[24]}) | (mul_22_8_n_29 & {in1[24]}));
 assign mul_22_8_n_307 = ~((mul_22_8_n_43 & {in2[11]}) | (mul_22_8_n_33 & {in1[12]}));
 assign mul_22_8_n_306 = ~((mul_22_8_n_45 & {in2[9]}) | (mul_22_8_n_32 & {in1[19]}));
 assign mul_22_8_n_305 = ~((mul_22_8_n_26 & {in2[9]}) | (mul_22_8_n_32 & {in1[18]}));
 assign mul_22_8_n_304 = ~((mul_22_8_n_26 & {in2[11]}) | (mul_22_8_n_33 & {in1[18]}));
 assign mul_22_8_n_303 = ~((mul_22_8_n_45 & {in2[11]}) | (mul_22_8_n_33 & {in1[19]}));
 assign mul_22_8_n_302 = ~(({in2[3]} & ~{in1[25]}) | (mul_22_8_n_29 & {in1[25]}));
 assign mul_22_8_n_301 = ~(({in2[5]} & ~{in1[26]}) | (mul_22_8_n_30 & {in1[26]}));
 assign mul_22_8_n_300 = ~((mul_22_8_n_26 & {in2[13]}) | (mul_22_8_n_10 & {in1[18]}));
 assign mul_22_8_n_298 = ~(({in1[16]} | mul_22_8_n_8) & ({in2[1]} | mul_22_8_n_24));
 assign mul_22_8_n_297 = ~((mul_22_8_n_23 & {in2[1]}) | (mul_22_8_n_8 & {in1[17]}));
 assign mul_22_8_n_296 = ~((mul_22_8_n_23 & {in2[3]}) | (mul_22_8_n_29 & {in1[17]}));
 assign mul_22_8_n_295 = ~((mul_22_8_n_24 & {in2[3]}) | (mul_22_8_n_29 & {in1[16]}));
 assign mul_22_8_n_294 = ~((mul_22_8_n_23 & {in2[5]}) | (mul_22_8_n_30 & {in1[17]}));
 assign mul_22_8_n_293 = ~((mul_22_8_n_24 & {in2[5]}) | (mul_22_8_n_30 & {in1[16]}));
 assign mul_22_8_n_292 = ~((mul_22_8_n_20 & {in2[11]}) | (mul_22_8_n_33 & {in1[13]}));
 assign mul_22_8_n_291 = ~((mul_22_8_n_23 & {in2[7]}) | (mul_22_8_n_31 & {in1[17]}));
 assign mul_22_8_n_290 = ~((mul_22_8_n_24 & {in2[7]}) | (mul_22_8_n_31 & {in1[16]}));
 assign mul_22_8_n_289 = ~((mul_22_8_n_24 & {in2[9]}) | (mul_22_8_n_32 & {in1[16]}));
 assign mul_22_8_n_288 = ~((mul_22_8_n_23 & {in2[9]}) | (mul_22_8_n_32 & {in1[17]}));
 assign mul_22_8_n_287 = ~((mul_22_8_n_24 & {in2[11]}) | (mul_22_8_n_33 & {in1[16]}));
 assign mul_22_8_n_286 = ~((mul_22_8_n_23 & {in2[11]}) | (mul_22_8_n_33 & {in1[17]}));
 assign mul_22_8_n_284 = ~(({in1[15]} | mul_22_8_n_8) & ({in2[1]} | mul_22_8_n_44));
 assign mul_22_8_n_283 = ~(({in1[14]} | mul_22_8_n_8) & ({in2[1]} | mul_22_8_n_22));
 assign mul_22_8_n_282 = ~((mul_22_8_n_24 & {in2[13]}) | (mul_22_8_n_10 & {in1[16]}));
 assign mul_22_8_n_281 = ~((mul_22_8_n_23 & {in2[13]}) | (mul_22_8_n_10 & {in1[17]}));
 assign mul_22_8_n_280 = ~((mul_22_8_n_44 & {in2[3]}) | (mul_22_8_n_29 & {in1[15]}));
 assign mul_22_8_n_279 = ~((mul_22_8_n_22 & {in2[3]}) | (mul_22_8_n_29 & {in1[14]}));
 assign mul_22_8_n_278 = ~((mul_22_8_n_44 & {in2[5]}) | (mul_22_8_n_30 & {in1[15]}));
 assign mul_22_8_n_277 = ~((mul_22_8_n_22 & {in2[5]}) | (mul_22_8_n_30 & {in1[14]}));
 assign mul_22_8_n_276 = ~(({in2[5]} & ~{in1[24]}) | (mul_22_8_n_30 & {in1[24]}));
 assign mul_22_8_n_275 = ~((mul_22_8_n_24 & {in2[15]}) | (mul_22_8_n_11 & {in1[16]}));
 assign mul_22_8_n_274 = ~((mul_22_8_n_22 & {in2[7]}) | (mul_22_8_n_31 & {in1[14]}));
 assign mul_22_8_n_273 = ~((mul_22_8_n_44 & {in2[7]}) | (mul_22_8_n_31 & {in1[15]}));
 assign mul_22_8_n_272 = ~((mul_22_8_n_22 & {in2[9]}) | (mul_22_8_n_32 & {in1[14]}));
 assign mul_22_8_n_271 = ~((mul_22_8_n_44 & {in2[9]}) | (mul_22_8_n_32 & {in1[15]}));
 assign mul_22_8_n_270 = ~(({in2[5]} & ~{in1[22]}) | (mul_22_8_n_30 & {in1[22]}));
 assign mul_22_8_n_269 = ~(({in1[12]} | mul_22_8_n_8) & ({in2[1]} | mul_22_8_n_43));
 assign mul_22_8_n_268 = ~(({in1[13]} | mul_22_8_n_8) & ({in2[1]} | mul_22_8_n_20));
 assign mul_22_8_n_267 = ~((mul_22_8_n_22 & {in2[11]}) | (mul_22_8_n_33 & {in1[14]}));
 assign mul_22_8_n_266 = ~((mul_22_8_n_44 & {in2[11]}) | (mul_22_8_n_33 & {in1[15]}));
 assign mul_22_8_n_265 = ~((mul_22_8_n_20 & {in2[3]}) | (mul_22_8_n_29 & {in1[13]}));
 assign mul_22_8_n_264 = ~((mul_22_8_n_43 & {in2[3]}) | (mul_22_8_n_29 & {in1[12]}));
 assign mul_22_8_n_263 = ~((mul_22_8_n_35 & {in2[29]}) | (mul_22_8_n_25 & {in1[1]}));
 assign mul_22_8_n_262 = ~((mul_22_8_n_19 & {in2[3]}) | (mul_22_8_n_29 & {in1[10]}));
 assign mul_22_8_n_261 = ~((mul_22_8_n_43 & {in2[5]}) | (mul_22_8_n_30 & {in1[12]}));
 assign mul_22_8_n_260 = ~((mul_22_8_n_20 & {in2[5]}) | (mul_22_8_n_30 & {in1[13]}));
 assign mul_22_8_n_259 = ~((mul_22_8_n_22 & {in2[13]}) | (mul_22_8_n_10 & {in1[14]}));
 assign mul_22_8_n_258 = ~((mul_22_8_n_44 & {in2[13]}) | (mul_22_8_n_10 & {in1[15]}));
 assign mul_22_8_n_257 = ~((mul_22_8_n_20 & {in2[7]}) | (mul_22_8_n_31 & {in1[13]}));
 assign mul_22_8_n_256 = ~((mul_22_8_n_43 & {in2[7]}) | (mul_22_8_n_31 & {in1[12]}));
 assign mul_22_8_n_255 = ~(({in2[1]} & ~{in1[25]}) | (mul_22_8_n_8 & {in1[25]}));
 assign mul_22_8_n_254 = ~((mul_22_8_n_15 & {in2[29]}) | (mul_22_8_n_25 & {in1[2]}));
 assign mul_22_8_n_253 = ~((mul_22_8_n_22 & {in2[15]}) | (mul_22_8_n_11 & {in1[14]}));
 assign mul_22_8_n_252 = ~((mul_22_8_n_44 & {in2[15]}) | (mul_22_8_n_11 & {in1[15]}));
 assign mul_22_8_n_251 = ~((mul_22_8_n_20 & {in2[9]}) | (mul_22_8_n_32 & {in1[13]}));
 assign mul_22_8_n_250 = ~((mul_22_8_n_43 & {in2[9]}) | (mul_22_8_n_32 & {in1[12]}));
 assign mul_22_8_n_249 = ~((mul_22_8_n_19 & {in2[1]}) | (mul_22_8_n_8 & {in1[10]}));
 assign mul_22_8_n_247 = ~(({in1[11]} | mul_22_8_n_8) & ({in2[1]} | mul_22_8_n_42));
 assign mul_22_8_n_246 = ~((mul_22_8_n_42 & {in2[3]}) | (mul_22_8_n_29 & {in1[11]}));
 assign mul_22_8_n_245 = ~((mul_22_8_n_25 & ~{in2[30]}) | ({in2[29]} & {in2[30]}));
 assign mul_22_8_n_244 = ~(({in2[27]} & ~{in2[28]}) | (mul_22_8_n_21 & {in2[28]}));
 assign mul_22_8_n_242 = ((mul_22_8_n_36 & ~{in2[22]}) | ({in2[21]} & {in2[22]}));
 assign mul_22_8_n_241 = ((mul_22_8_n_13 & ~{in2[20]}) | ({in2[19]} & {in2[20]}));
 assign mul_22_8_n_240 = ((mul_22_8_n_12 & ~{in2[18]}) | ({in2[17]} & {in2[18]}));
 assign mul_22_8_n_239 = ((mul_22_8_n_11 & ~{in2[16]}) | ({in2[15]} & {in2[16]}));
 assign mul_22_8_n_238 = ((mul_22_8_n_10 & ~{in2[14]}) | ({in2[13]} & {in2[14]}));
 assign mul_22_8_n_237 = ((mul_22_8_n_33 & ~{in2[12]}) | ({in2[11]} & {in2[12]}));
 assign mul_22_8_n_236 = ((mul_22_8_n_32 & ~{in2[10]}) | ({in2[9]} & {in2[10]}));
 assign mul_22_8_n_235 = ((mul_22_8_n_31 & ~{in2[8]}) | ({in2[7]} & {in2[8]}));
 assign mul_22_8_n_234 = ((mul_22_8_n_30 & ~{in2[6]}) | ({in2[5]} & {in2[6]}));
 assign mul_22_8_n_233 = ((mul_22_8_n_29 & ~{in2[4]}) | ({in2[3]} & {in2[4]}));
 assign mul_22_8_n_232 = ((mul_22_8_n_8 & ~{in2[2]}) | ({in2[1]} & {in2[2]}));
 assign mul_22_8_n_196 = ~mul_22_8_n_195;
 assign mul_22_8_n_87 = ~mul_22_8_n_86;
 assign mul_22_8_n_73 = ~mul_22_8_n_72;
 assign mul_22_8_n_71 = ~mul_22_8_n_70;
 assign mul_22_8_n_69 = ~((mul_22_8_n_38 & {in2[25]}) | (mul_22_8_n_18 & {in1[7]}));
 assign mul_22_8_n_68 = ~((mul_22_8_n_9 & {in2[23]}) | (mul_22_8_n_17 & {in1[0]}));
 assign mul_22_8_n_67 = ~((mul_22_8_n_37 & {in2[27]}) | (mul_22_8_n_21 & {in1[5]}));
 assign mul_22_8_n_66 = ~((mul_22_8_n_9 & {in2[21]}) | (mul_22_8_n_36 & {in1[0]}));
 assign mul_22_8_n_64 = ~((mul_22_8_n_42 & {in2[21]}) | (mul_22_8_n_36 & {in1[11]}));
 assign mul_22_8_n_63 = ~((mul_22_8_n_9 & {in2[19]}) | (mul_22_8_n_13 & {in1[0]}));
 assign mul_22_8_n_62 = ~((mul_22_8_n_9 & {in2[17]}) | (mul_22_8_n_12 & {in1[0]}));
 assign mul_22_8_n_61 = ~((mul_22_8_n_9 & {in2[15]}) | (mul_22_8_n_11 & {in1[0]}));
 assign mul_22_8_n_60 = ~((mul_22_8_n_20 & {in2[19]}) | (mul_22_8_n_13 & {in1[13]}));
 assign mul_22_8_n_59 = ~((mul_22_8_n_40 & {in2[23]}) | (mul_22_8_n_17 & {in1[9]}));
 assign mul_22_8_n_58 = ~((mul_22_8_n_9 & {in2[13]}) | (mul_22_8_n_10 & {in1[0]}));
 assign mul_22_8_n_57 = ~((mul_22_8_n_9 & {in2[11]}) | (mul_22_8_n_33 & {in1[0]}));
 assign mul_22_8_n_56 = ~((mul_22_8_n_9 & {in2[9]}) | (mul_22_8_n_32 & {in1[0]}));
 assign mul_22_8_n_55 = ~(({in1[0]} | mul_22_8_n_8) & ({in2[1]} | mul_22_8_n_9));
 assign mul_22_8_n_54 = ~((mul_22_8_n_9 & {in2[7]}) | (mul_22_8_n_31 & {in1[0]}));
 assign mul_22_8_n_53 = ~((mul_22_8_n_9 & {in2[3]}) | (mul_22_8_n_29 & {in1[0]}));
 assign mul_22_8_n_52 = ~((mul_22_8_n_9 & {in2[5]}) | (mul_22_8_n_30 & {in1[0]}));
 assign mul_22_8_n_51 = ~({in2[30]} ^ {in2[31]});
 assign mul_22_8_n_205 = ~((mul_22_8_n_40 & {in2[9]}) | (mul_22_8_n_32 & {in1[9]}));
 assign mul_22_8_n_204 = ~((mul_22_8_n_41 & {in2[9]}) | (mul_22_8_n_32 & {in1[8]}));
 assign mul_22_8_n_203 = ~((mul_22_8_n_39 & {in2[5]}) | (mul_22_8_n_30 & {in1[6]}));
 assign mul_22_8_n_202 = ~((mul_22_8_n_38 & {in2[5]}) | (mul_22_8_n_30 & {in1[7]}));
 assign mul_22_8_n_201 = ~((mul_22_8_n_19 & {in2[15]}) | (mul_22_8_n_11 & {in1[10]}));
 assign mul_22_8_n_200 = ~((mul_22_8_n_42 & {in2[15]}) | (mul_22_8_n_11 & {in1[11]}));
 assign mul_22_8_n_199 = ~((mul_22_8_n_40 & {in2[11]}) | (mul_22_8_n_33 & {in1[9]}));
 assign mul_22_8_n_198 = ~((mul_22_8_n_41 & {in2[11]}) | (mul_22_8_n_33 & {in1[8]}));
 assign mul_22_8_n_197 = ~(({in1[5]} | mul_22_8_n_8) & ({in2[1]} | mul_22_8_n_37));
 assign mul_22_8_n_195 = ~(({in1[4]} | mul_22_8_n_8) & ({in2[1]} | mul_22_8_n_16));
 assign mul_22_8_n_194 = ~((mul_22_8_n_35 & {in2[27]}) | (mul_22_8_n_21 & {in1[1]}));
 assign mul_22_8_n_193 = ~((mul_22_8_n_39 & {in2[7]}) | (mul_22_8_n_31 & {in1[6]}));
 assign mul_22_8_n_192 = ~((mul_22_8_n_38 & {in2[7]}) | (mul_22_8_n_31 & {in1[7]}));
 assign mul_22_8_n_191 = ~((mul_22_8_n_16 & {in2[11]}) | (mul_22_8_n_33 & {in1[4]}));
 assign mul_22_8_n_190 = ~((mul_22_8_n_43 & {in2[19]}) | (mul_22_8_n_13 & {in1[12]}));
 assign mul_22_8_n_189 = ~((mul_22_8_n_41 & {in2[3]}) | (mul_22_8_n_29 & {in1[8]}));
 assign mul_22_8_n_188 = ~((mul_22_8_n_16 & {in2[3]}) | (mul_22_8_n_29 & {in1[4]}));
 assign mul_22_8_n_187 = ~((mul_22_8_n_37 & {in2[3]}) | (mul_22_8_n_29 & {in1[5]}));
 assign mul_22_8_n_186 = ~((mul_22_8_n_40 & {in2[13]}) | (mul_22_8_n_10 & {in1[9]}));
 assign mul_22_8_n_185 = ~((mul_22_8_n_41 & {in2[13]}) | (mul_22_8_n_10 & {in1[8]}));
 assign mul_22_8_n_184 = ~((mul_22_8_n_39 & {in2[9]}) | (mul_22_8_n_32 & {in1[6]}));
 assign mul_22_8_n_183 = ~((mul_22_8_n_38 & {in2[9]}) | (mul_22_8_n_32 & {in1[7]}));
 assign mul_22_8_n_182 = ~((mul_22_8_n_42 & {in2[17]}) | (mul_22_8_n_12 & {in1[11]}));
 assign mul_22_8_n_181 = ~((mul_22_8_n_19 & {in2[17]}) | (mul_22_8_n_12 & {in1[10]}));
 assign mul_22_8_n_180 = ~((mul_22_8_n_37 & {in2[5]}) | (mul_22_8_n_30 & {in1[5]}));
 assign mul_22_8_n_179 = ~((mul_22_8_n_16 & {in2[5]}) | (mul_22_8_n_30 & {in1[4]}));
 assign mul_22_8_n_178 = ~((mul_22_8_n_15 & {in2[27]}) | (mul_22_8_n_21 & {in1[2]}));
 assign mul_22_8_n_177 = ~((mul_22_8_n_14 & {in2[27]}) | (mul_22_8_n_21 & {in1[3]}));
 assign mul_22_8_n_176 = ~(({in1[2]} | mul_22_8_n_8) & ({in2[1]} | mul_22_8_n_15));
 assign mul_22_8_n_175 = ~((mul_22_8_n_14 & {in2[1]}) | (mul_22_8_n_8 & {in1[3]}));
 assign mul_22_8_n_174 = ~((mul_22_8_n_38 & {in2[11]}) | (mul_22_8_n_33 & {in1[7]}));
 assign mul_22_8_n_173 = ~((mul_22_8_n_39 & {in2[11]}) | (mul_22_8_n_33 & {in1[6]}));
 assign mul_22_8_n_172 = ~((mul_22_8_n_37 & {in2[7]}) | (mul_22_8_n_31 & {in1[5]}));
 assign mul_22_8_n_171 = ~((mul_22_8_n_16 & {in2[7]}) | (mul_22_8_n_31 & {in1[4]}));
 assign mul_22_8_n_170 = ~((mul_22_8_n_41 & {in2[15]}) | (mul_22_8_n_11 & {in1[8]}));
 assign mul_22_8_n_169 = ~((mul_22_8_n_40 & {in2[15]}) | (mul_22_8_n_11 & {in1[9]}));
 assign mul_22_8_n_168 = ~((mul_22_8_n_14 & {in2[3]}) | (mul_22_8_n_29 & {in1[3]}));
 assign mul_22_8_n_167 = ~((mul_22_8_n_15 & {in2[3]}) | (mul_22_8_n_29 & {in1[2]}));
 assign mul_22_8_n_166 = ~((mul_22_8_n_16 & {in2[27]}) | (mul_22_8_n_21 & {in1[4]}));
 assign mul_22_8_n_165 = ~((mul_22_8_n_40 & {in2[3]}) | (mul_22_8_n_29 & {in1[9]}));
 assign mul_22_8_n_164 = ~((mul_22_8_n_16 & {in2[9]}) | (mul_22_8_n_32 & {in1[4]}));
 assign mul_22_8_n_163 = ~((mul_22_8_n_37 & {in2[9]}) | (mul_22_8_n_32 & {in1[5]}));
 assign mul_22_8_n_162 = ~((mul_22_8_n_15 & {in2[5]}) | (mul_22_8_n_30 & {in1[2]}));
 assign mul_22_8_n_161 = ~((mul_22_8_n_14 & {in2[5]}) | (mul_22_8_n_30 & {in1[3]}));
 assign mul_22_8_n_160 = ~((mul_22_8_n_38 & {in2[13]}) | (mul_22_8_n_10 & {in1[7]}));
 assign mul_22_8_n_159 = ~((mul_22_8_n_39 & {in2[13]}) | (mul_22_8_n_10 & {in1[6]}));
 assign mul_22_8_n_158 = ~(({in1[1]} | mul_22_8_n_8) & ({in2[1]} | mul_22_8_n_35));
 assign mul_22_8_n_157 = ~((mul_22_8_n_19 & {in2[19]}) | (mul_22_8_n_13 & {in1[10]}));
 assign mul_22_8_n_156 = ~((mul_22_8_n_42 & {in2[19]}) | (mul_22_8_n_13 & {in1[11]}));
 assign mul_22_8_n_155 = ~((mul_22_8_n_14 & {in2[7]}) | (mul_22_8_n_31 & {in1[3]}));
 assign mul_22_8_n_154 = ~((mul_22_8_n_15 & {in2[7]}) | (mul_22_8_n_31 & {in1[2]}));
 assign mul_22_8_n_153 = ~((mul_22_8_n_43 & {in2[15]}) | (mul_22_8_n_11 & {in1[12]}));
 assign mul_22_8_n_152 = ~((mul_22_8_n_35 & {in2[3]}) | (mul_22_8_n_29 & {in1[1]}));
 assign mul_22_8_n_151 = ~((mul_22_8_n_41 & {in2[17]}) | (mul_22_8_n_12 & {in1[8]}));
 assign mul_22_8_n_150 = ~((mul_22_8_n_40 & {in2[17]}) | (mul_22_8_n_12 & {in1[9]}));
 assign mul_22_8_n_149 = ~((mul_22_8_n_37 & {in2[11]}) | (mul_22_8_n_33 & {in1[5]}));
 assign mul_22_8_n_148 = ~((mul_22_8_n_19 & {in2[9]}) | (mul_22_8_n_32 & {in1[10]}));
 assign mul_22_8_n_147 = ~((mul_22_8_n_35 & {in2[5]}) | (mul_22_8_n_30 & {in1[1]}));
 assign mul_22_8_n_146 = ~((mul_22_8_n_39 & {in2[15]}) | (mul_22_8_n_11 & {in1[6]}));
 assign mul_22_8_n_145 = ~((mul_22_8_n_38 & {in2[15]}) | (mul_22_8_n_11 & {in1[7]}));
 assign mul_22_8_n_144 = ~((mul_22_8_n_15 & {in2[9]}) | (mul_22_8_n_32 & {in1[2]}));
 assign mul_22_8_n_143 = ~((mul_22_8_n_14 & {in2[9]}) | (mul_22_8_n_32 & {in1[3]}));
 assign mul_22_8_n_142 = ~((mul_22_8_n_37 & {in2[13]}) | (mul_22_8_n_10 & {in1[5]}));
 assign mul_22_8_n_141 = ~((mul_22_8_n_16 & {in2[13]}) | (mul_22_8_n_10 & {in1[4]}));
 assign mul_22_8_n_140 = ~((mul_22_8_n_20 & {in2[15]}) | (mul_22_8_n_11 & {in1[13]}));
 assign mul_22_8_n_139 = ~((mul_22_8_n_35 & {in2[7]}) | (mul_22_8_n_31 & {in1[1]}));
 assign mul_22_8_n_138 = ~((mul_22_8_n_19 & {in2[21]}) | (mul_22_8_n_36 & {in1[10]}));
 assign mul_22_8_n_137 = ~((mul_22_8_n_40 & {in2[5]}) | (mul_22_8_n_30 & {in1[9]}));
 assign mul_22_8_n_136 = ~((mul_22_8_n_15 & {in2[11]}) | (mul_22_8_n_33 & {in1[2]}));
 assign mul_22_8_n_135 = ~((mul_22_8_n_14 & {in2[11]}) | (mul_22_8_n_33 & {in1[3]}));
 assign mul_22_8_n_134 = ~((mul_22_8_n_41 & {in2[19]}) | (mul_22_8_n_13 & {in1[8]}));
 assign mul_22_8_n_133 = ~((mul_22_8_n_40 & {in2[19]}) | (mul_22_8_n_13 & {in1[9]}));
 assign mul_22_8_n_132 = ~((mul_22_8_n_38 & {in2[17]}) | (mul_22_8_n_12 & {in1[7]}));
 assign mul_22_8_n_131 = ~((mul_22_8_n_39 & {in2[17]}) | (mul_22_8_n_12 & {in1[6]}));
 assign mul_22_8_n_130 = ~((mul_22_8_n_35 & {in2[9]}) | (mul_22_8_n_32 & {in1[1]}));
 assign mul_22_8_n_129 = ~((mul_22_8_n_35 & {in2[25]}) | (mul_22_8_n_18 & {in1[1]}));
 assign mul_22_8_n_128 = ~((mul_22_8_n_41 & {in2[5]}) | (mul_22_8_n_30 & {in1[8]}));
 assign mul_22_8_n_127 = ~((mul_22_8_n_37 & {in2[15]}) | (mul_22_8_n_11 & {in1[5]}));
 assign mul_22_8_n_126 = ~((mul_22_8_n_16 & {in2[15]}) | (mul_22_8_n_11 & {in1[4]}));
 assign mul_22_8_n_125 = ~((mul_22_8_n_14 & {in2[13]}) | (mul_22_8_n_10 & {in1[3]}));
 assign mul_22_8_n_124 = ~((mul_22_8_n_15 & {in2[13]}) | (mul_22_8_n_10 & {in1[2]}));
 assign mul_22_8_n_123 = ~((mul_22_8_n_35 & {in2[11]}) | (mul_22_8_n_33 & {in1[1]}));
 assign mul_22_8_n_122 = ~((mul_22_8_n_15 & {in2[25]}) | (mul_22_8_n_18 & {in1[2]}));
 assign mul_22_8_n_121 = ~((mul_22_8_n_14 & {in2[25]}) | (mul_22_8_n_18 & {in1[3]}));
 assign mul_22_8_n_120 = ~((mul_22_8_n_39 & {in2[19]}) | (mul_22_8_n_13 & {in1[6]}));
 assign mul_22_8_n_119 = ~((mul_22_8_n_38 & {in2[19]}) | (mul_22_8_n_13 & {in1[7]}));
 assign mul_22_8_n_118 = ~((mul_22_8_n_37 & {in2[17]}) | (mul_22_8_n_12 & {in1[5]}));
 assign mul_22_8_n_117 = ~((mul_22_8_n_16 & {in2[17]}) | (mul_22_8_n_12 & {in1[4]}));
 assign mul_22_8_n_116 = ~((mul_22_8_n_15 & {in2[15]}) | (mul_22_8_n_11 & {in1[2]}));
 assign mul_22_8_n_115 = ~((mul_22_8_n_14 & {in2[15]}) | (mul_22_8_n_11 & {in1[3]}));
 assign mul_22_8_n_114 = ~((mul_22_8_n_40 & {in2[21]}) | (mul_22_8_n_36 & {in1[9]}));
 assign mul_22_8_n_113 = ~((mul_22_8_n_41 & {in2[21]}) | (mul_22_8_n_36 & {in1[8]}));
 assign mul_22_8_n_112 = ~((mul_22_8_n_35 & {in2[13]}) | (mul_22_8_n_10 & {in1[1]}));
 assign mul_22_8_n_111 = ~((mul_22_8_n_19 & {in2[11]}) | (mul_22_8_n_33 & {in1[10]}));
 assign mul_22_8_n_110 = ~((mul_22_8_n_37 & {in2[25]}) | (mul_22_8_n_18 & {in1[5]}));
 assign mul_22_8_n_109 = ~((mul_22_8_n_16 & {in2[25]}) | (mul_22_8_n_18 & {in1[4]}));
 assign mul_22_8_n_108 = ~((mul_22_8_n_35 & {in2[15]}) | (mul_22_8_n_11 & {in1[1]}));
 assign mul_22_8_n_107 = ~((mul_22_8_n_15 & {in2[17]}) | (mul_22_8_n_12 & {in1[2]}));
 assign mul_22_8_n_106 = ~((mul_22_8_n_14 & {in2[17]}) | (mul_22_8_n_12 & {in1[3]}));
 assign mul_22_8_n_105 = ~((mul_22_8_n_37 & {in2[19]}) | (mul_22_8_n_13 & {in1[5]}));
 assign mul_22_8_n_104 = ~((mul_22_8_n_16 & {in2[19]}) | (mul_22_8_n_13 & {in1[4]}));
 assign mul_22_8_n_103 = ~((mul_22_8_n_42 & {in2[11]}) | (mul_22_8_n_33 & {in1[11]}));
 assign mul_22_8_n_102 = ~((mul_22_8_n_38 & {in2[21]}) | (mul_22_8_n_36 & {in1[7]}));
 assign mul_22_8_n_101 = ~((mul_22_8_n_39 & {in2[21]}) | (mul_22_8_n_36 & {in1[6]}));
 assign mul_22_8_n_100 = ~((mul_22_8_n_35 & {in2[23]}) | (mul_22_8_n_17 & {in1[1]}));
 assign mul_22_8_n_99 = ~((mul_22_8_n_40 & {in2[7]}) | (mul_22_8_n_31 & {in1[9]}));
 assign mul_22_8_n_98 = ~((mul_22_8_n_39 & {in2[25]}) | (mul_22_8_n_18 & {in1[6]}));
 assign mul_22_8_n_97 = ~((mul_22_8_n_41 & {in2[23]}) | (mul_22_8_n_17 & {in1[8]}));
 assign mul_22_8_n_96 = ~((mul_22_8_n_41 & {in2[7]}) | (mul_22_8_n_31 & {in1[8]}));
 assign mul_22_8_n_95 = ~((mul_22_8_n_35 & {in2[17]}) | (mul_22_8_n_12 & {in1[1]}));
 assign mul_22_8_n_94 = ~((mul_22_8_n_15 & {in2[19]}) | (mul_22_8_n_13 & {in1[2]}));
 assign mul_22_8_n_93 = ~((mul_22_8_n_14 & {in2[19]}) | (mul_22_8_n_13 & {in1[3]}));
 assign mul_22_8_n_92 = ~(({in1[6]} | mul_22_8_n_8) & ({in2[1]} | mul_22_8_n_39));
 assign mul_22_8_n_91 = ~((mul_22_8_n_14 & {in2[23]}) | (mul_22_8_n_17 & {in1[3]}));
 assign mul_22_8_n_90 = ~((mul_22_8_n_15 & {in2[23]}) | (mul_22_8_n_17 & {in1[2]}));
 assign mul_22_8_n_89 = ~((mul_22_8_n_37 & {in2[21]}) | (mul_22_8_n_36 & {in1[5]}));
 assign mul_22_8_n_88 = ~((mul_22_8_n_16 & {in2[21]}) | (mul_22_8_n_36 & {in1[4]}));
 assign mul_22_8_n_86 = ~((mul_22_8_n_38 & {in2[1]}) | (mul_22_8_n_8 & {in1[7]}));
 assign mul_22_8_n_85 = ~((mul_22_8_n_35 & {in2[19]}) | (mul_22_8_n_13 & {in1[1]}));
 assign mul_22_8_n_84 = ~((mul_22_8_n_38 & {in2[23]}) | (mul_22_8_n_17 & {in1[7]}));
 assign mul_22_8_n_83 = ~((mul_22_8_n_39 & {in2[23]}) | (mul_22_8_n_17 & {in1[6]}));
 assign mul_22_8_n_82 = ~((mul_22_8_n_16 & {in2[23]}) | (mul_22_8_n_17 & {in1[4]}));
 assign mul_22_8_n_81 = ~((mul_22_8_n_37 & {in2[23]}) | (mul_22_8_n_17 & {in1[5]}));
 assign mul_22_8_n_80 = ~((mul_22_8_n_15 & {in2[21]}) | (mul_22_8_n_36 & {in1[2]}));
 assign mul_22_8_n_79 = ~((mul_22_8_n_14 & {in2[21]}) | (mul_22_8_n_36 & {in1[3]}));
 assign mul_22_8_n_78 = ~((mul_22_8_n_43 & {in2[17]}) | (mul_22_8_n_12 & {in1[12]}));
 assign mul_22_8_n_77 = ~((mul_22_8_n_35 & {in2[21]}) | (mul_22_8_n_36 & {in1[1]}));
 assign mul_22_8_n_76 = ~((mul_22_8_n_20 & {in2[17]}) | (mul_22_8_n_12 & {in1[13]}));
 assign mul_22_8_n_75 = ~((mul_22_8_n_19 & {in2[13]}) | (mul_22_8_n_10 & {in1[10]}));
 assign mul_22_8_n_74 = ~((mul_22_8_n_42 & {in2[13]}) | (mul_22_8_n_10 & {in1[11]}));
 assign mul_22_8_n_72 = ~(({in1[6]} | mul_22_8_n_29) & ({in2[3]} | mul_22_8_n_39));
 assign mul_22_8_n_70 = ~((mul_22_8_n_38 & {in2[3]}) | (mul_22_8_n_29 & {in1[7]}));
 assign mul_22_8_n_50 = ~({in2[26]} | mul_22_8_n_21);
 assign mul_22_8_n_49 = ~({in2[28]} | mul_22_8_n_25);
 assign mul_22_8_n_48 = ~({in2[31]} | mul_22_8_n_35);
 assign asc001_0_ = ~(mul_22_8_n_34 | mul_22_8_n_9);
 assign mul_22_8_n_46 = ~{in1[20]};
 assign mul_22_8_n_45 = ~{in1[19]};
 assign mul_22_8_n_44 = ~{in1[15]};
 assign mul_22_8_n_43 = ~{in1[12]};
 assign mul_22_8_n_42 = ~{in1[11]};
 assign mul_22_8_n_41 = ~{in1[8]};
 assign mul_22_8_n_40 = ~{in1[9]};
 assign mul_22_8_n_39 = ~{in1[6]};
 assign mul_22_8_n_38 = ~{in1[7]};
 assign mul_22_8_n_37 = ~{in1[5]};
 assign mul_22_8_n_36 = ~{in2[21]};
 assign mul_22_8_n_35 = ~{in1[1]};
 assign mul_22_8_n_34 = ~{in2[0]};
 assign mul_22_8_n_33 = ~{in2[11]};
 assign mul_22_8_n_32 = ~{in2[9]};
 assign mul_22_8_n_31 = ~{in2[7]};
 assign mul_22_8_n_30 = ~{in2[5]};
 assign mul_22_8_n_29 = ~{in2[3]};
 assign mul_22_8_n_27 = ~{in1[21]};
 assign mul_22_8_n_26 = ~{in1[18]};
 assign mul_22_8_n_25 = ~{in2[29]};
 assign mul_22_8_n_24 = ~{in1[16]};
 assign mul_22_8_n_23 = ~{in1[17]};
 assign mul_22_8_n_22 = ~{in1[14]};
 assign mul_22_8_n_21 = ~{in2[27]};
 assign mul_22_8_n_20 = ~{in1[13]};
 assign mul_22_8_n_19 = ~{in1[10]};
 assign mul_22_8_n_18 = ~{in2[25]};
 assign mul_22_8_n_17 = ~{in2[23]};
 assign mul_22_8_n_16 = ~{in1[4]};
 assign mul_22_8_n_15 = ~{in1[2]};
 assign mul_22_8_n_14 = ~{in1[3]};
 assign mul_22_8_n_13 = ~{in2[19]};
 assign mul_22_8_n_12 = ~{in2[17]};
 assign mul_22_8_n_11 = ~{in2[15]};
 assign mul_22_8_n_10 = ~{in2[13]};
 assign mul_22_8_n_9 = ~{in1[0]};
 assign mul_22_8_n_8 = ~{in2[1]};
 assign mul_22_8_n_6 = (mul_22_8_n_837 | mul_22_8_n_839);
 assign mul_22_8_n_5 = (n_38 | n_28);
 assign mul_22_8_n_4 = (n_36 | n_81);
 assign asc001_16_ = (mul_22_8_n_808 ^ mul_22_8_n_827);
 assign mul_22_8_n_2 = (mul_22_8_n_1280 & mul_22_8_n_1304);
 assign mul_22_8_n_1 = ~(n_65 & (~n_86 | n_67));
 assign mul_22_8_n_0 = ~(({in2[25]} & ~{in2[26]}) | (mul_22_8_n_18 & {in2[26]}));
 assign n_0 = ~clr;
 assign n_154 = ~(mul_22_8_n_887 & (mul_22_8_n_885 | (mul_22_8_n_898 & mul_22_8_n_886)));
 assign n_155 = ~(({in2[23]} & ~{in2[24]}) | (mul_22_8_n_17 & {in2[24]}));
 assign mul_22_8_n_939 = (mul_22_8_n_636 ^ (mul_22_8_n_631 ^ mul_22_8_n_639));
 assign mul_22_8_n_938 = (mul_22_8_n_646 ^ (mul_22_8_n_643 ^ mul_22_8_n_645));
 assign mul_22_8_n_937 = (mul_22_8_n_642 ^ (mul_22_8_n_635 ^ mul_22_8_n_638));
 assign mul_22_8_n_936 = (mul_22_8_n_644 ^ (mul_22_8_n_629 ^ mul_22_8_n_633));
 assign mul_22_8_n_935 = (mul_22_8_n_625 ^ (mul_22_8_n_624 ^ mul_22_8_n_641));
 assign mul_22_8_n_1292 = (n_25 ^ (n_51 ^ n_68));
 assign mul_22_8_n_932 = (mul_22_8_n_940 ^ (mul_22_8_n_941 ^ mul_22_8_n_942));
 assign mul_22_8_n_931 = (mul_22_8_n_943 ^ (mul_22_8_n_944 ^ mul_22_8_n_707));
 assign mul_22_8_n_928 = (mul_22_8_n_937 ^ (mul_22_8_n_938 ^ mul_22_8_n_939));
 assign mul_22_8_n_924 = (mul_22_8_n_931 ^ (mul_22_8_n_932 ^ mul_22_8_n_933));
 assign mul_22_8_n_923 = (mul_22_8_n_928 ^ (mul_22_8_n_929 ^ mul_22_8_n_930));
 assign mul_22_8_n_927 = (mul_22_8_n_934 ^ (mul_22_8_n_935 ^ mul_22_8_n_936));
 assign mul_22_8_n_921 = (mul_22_8_n_925 ^ (mul_22_8_n_926 ^ mul_22_8_n_927));
 assign mul_22_8_n_920 = (mul_22_8_n_922 ^ (mul_22_8_n_923 ^ mul_22_8_n_924));
endmodule


