`timescale 1ps / 1ps
module vitdodec_Mod_32Ux32U_32U_4(
          in2,
          in1,
          out1,
          clk,
          clr
);
   input [31:0] in2;
   input [31:0] in1;
   output [31:0] out1;
   input clk;
   input clr;
wire sub_181_2_n_0, sub_181_2_n_22, sub_181_2_n_28, sub_181_2_n_29,
     sub_181_2_n_30, sub_200_2_n_0, sub_200_2_n_1, sub_200_2_n_2, sub_200_2_n_5,
     sub_200_2_n_6, sub_200_2_n_8, sub_200_2_n_16, sub_200_2_n_27,
     sub_200_2_n_28, sub_200_2_n_32, sub_200_2_n_33, sub_200_2_n_35,
     sub_200_2_n_36, sub_200_2_n_37, sub_219_2_n_3, sub_219_2_n_4, sub_219_2_n_5,
     sub_219_2_n_9, sub_219_2_n_17, sub_219_2_n_26, sub_219_2_n_29,
     sub_219_2_n_37, sub_219_2_n_38, sub_219_2_n_39, sub_219_2_n_41,
     sub_219_2_n_44, sub_238_2_n_0, sub_238_2_n_1, sub_238_2_n_2, sub_238_2_n_3,
     sub_238_2_n_4, sub_238_2_n_8, sub_238_2_n_9, sub_238_2_n_12, sub_238_2_n_14,
     sub_238_2_n_15, sub_238_2_n_16, sub_238_2_n_17, sub_238_2_n_19,
     sub_238_2_n_23, sub_238_2_n_24, sub_238_2_n_25, sub_238_2_n_26,
     sub_238_2_n_28, sub_238_2_n_30, sub_238_2_n_31, sub_238_2_n_33,
     sub_238_2_n_34, sub_238_2_n_36, sub_238_2_n_37, sub_238_2_n_38,
     sub_257_2_n_1, sub_257_2_n_2, sub_257_2_n_3, sub_257_2_n_4, sub_257_2_n_5,
     sub_257_2_n_6, sub_257_2_n_8, sub_257_2_n_9, sub_257_2_n_10, sub_257_2_n_11,
     sub_257_2_n_15, sub_257_2_n_16, sub_257_2_n_17, sub_257_2_n_18,
     sub_257_2_n_19, sub_257_2_n_22, sub_257_2_n_24, sub_257_2_n_25,
     sub_257_2_n_27, sub_257_2_n_31, sub_257_2_n_32, sub_257_2_n_33,
     sub_257_2_n_34, sub_257_2_n_35, sub_257_2_n_36, sub_257_2_n_37,
     sub_257_2_n_39, sub_257_2_n_41, sub_257_2_n_43, sub_257_2_n_44,
     sub_257_2_n_45, sub_257_2_n_48, sub_257_2_n_49, sub_276_2_n_0,
     sub_276_2_n_1, sub_276_2_n_2, sub_276_2_n_3, sub_276_2_n_4, sub_276_2_n_5,
     sub_276_2_n_6, sub_276_2_n_7, sub_276_2_n_9, sub_276_2_n_11, sub_276_2_n_12,
     sub_276_2_n_13, sub_276_2_n_16, sub_276_2_n_17, sub_276_2_n_18,
     sub_276_2_n_19, sub_276_2_n_23, sub_276_2_n_24, sub_276_2_n_25,
     sub_276_2_n_26, sub_276_2_n_27, sub_276_2_n_28, sub_276_2_n_35,
     sub_276_2_n_36, sub_276_2_n_37, sub_276_2_n_38, sub_276_2_n_40,
     sub_276_2_n_43, sub_276_2_n_47, sub_276_2_n_48, sub_276_2_n_50,
     sub_276_2_n_51, sub_276_2_n_52, sub_276_2_n_54, sub_276_2_n_55,
     sub_276_2_n_56, sub_295_2_n_0, sub_295_2_n_1, sub_295_2_n_2, sub_295_2_n_3,
     sub_295_2_n_4, sub_295_2_n_6, sub_295_2_n_7, sub_295_2_n_8, sub_295_2_n_9,
     sub_295_2_n_10, sub_295_2_n_13, sub_295_2_n_14, sub_295_2_n_15,
     sub_295_2_n_16, sub_295_2_n_19, sub_295_2_n_20, sub_295_2_n_21,
     sub_295_2_n_22, sub_295_2_n_23, sub_295_2_n_24, sub_295_2_n_25,
     sub_295_2_n_28, sub_295_2_n_29, sub_295_2_n_30, sub_295_2_n_31,
     sub_295_2_n_32, sub_295_2_n_33, sub_295_2_n_39, sub_295_2_n_40,
     sub_295_2_n_41, sub_295_2_n_43, sub_295_2_n_44, sub_295_2_n_45,
     sub_295_2_n_49, sub_295_2_n_51, sub_295_2_n_53, sub_295_2_n_54,
     sub_295_2_n_55, sub_295_2_n_57, sub_295_2_n_58, sub_295_2_n_59,
     sub_295_2_n_62, sub_314_2_n_0, sub_314_2_n_1, sub_314_2_n_2, sub_314_2_n_3,
     sub_314_2_n_4, sub_314_2_n_5, sub_314_2_n_6, sub_314_2_n_7, sub_314_2_n_8,
     sub_314_2_n_9, sub_314_2_n_10, sub_314_2_n_12, sub_314_2_n_13,
     sub_314_2_n_17, sub_314_2_n_18, sub_314_2_n_19, sub_314_2_n_20,
     sub_314_2_n_21, sub_314_2_n_22, sub_314_2_n_23, sub_314_2_n_24,
     sub_314_2_n_25, sub_314_2_n_27, sub_314_2_n_28, sub_314_2_n_29,
     sub_314_2_n_30, sub_314_2_n_31, sub_314_2_n_32, sub_314_2_n_33,
     sub_314_2_n_35, sub_314_2_n_37, sub_314_2_n_38, sub_314_2_n_39,
     sub_314_2_n_40, sub_314_2_n_41, sub_314_2_n_42, sub_314_2_n_44,
     sub_314_2_n_45, sub_314_2_n_48, sub_314_2_n_50, sub_314_2_n_52,
     sub_314_2_n_53, sub_314_2_n_55, sub_314_2_n_57, sub_314_2_n_58,
     sub_314_2_n_59, sub_314_2_n_60, sub_314_2_n_63, sub_314_2_n_64,
     sub_314_2_n_67, sub_314_2_n_68, sub_333_2_n_0, sub_333_2_n_1, sub_333_2_n_2,
     sub_333_2_n_3, sub_333_2_n_4, sub_333_2_n_5, sub_333_2_n_6, sub_333_2_n_7,
     sub_333_2_n_8, sub_333_2_n_9, sub_333_2_n_10, sub_333_2_n_11,
     sub_333_2_n_12, sub_333_2_n_14, sub_333_2_n_16, sub_333_2_n_18,
     sub_333_2_n_19, sub_333_2_n_20, sub_333_2_n_21, sub_333_2_n_22,
     sub_333_2_n_23, sub_333_2_n_24, sub_333_2_n_25, sub_333_2_n_27,
     sub_333_2_n_28, sub_333_2_n_29, sub_333_2_n_30, sub_333_2_n_31,
     sub_333_2_n_33, sub_333_2_n_34, sub_333_2_n_35, sub_333_2_n_37,
     sub_333_2_n_39, sub_333_2_n_41, sub_333_2_n_42, sub_333_2_n_43,
     sub_333_2_n_44, sub_333_2_n_46, sub_333_2_n_47, sub_333_2_n_48,
     sub_333_2_n_49, sub_333_2_n_52, sub_333_2_n_54, sub_333_2_n_55,
     sub_333_2_n_56, sub_333_2_n_58, sub_333_2_n_59, sub_333_2_n_60,
     sub_333_2_n_62, sub_333_2_n_63, sub_333_2_n_65, sub_333_2_n_67,
     sub_333_2_n_70, sub_333_2_n_75, sub_333_2_n_76, sub_333_2_n_78,
     sub_352_2_n_1, sub_352_2_n_2, sub_352_2_n_3, sub_352_2_n_4, sub_352_2_n_5,
     sub_352_2_n_6, sub_352_2_n_7, sub_352_2_n_8, sub_352_2_n_9, sub_352_2_n_10,
     sub_352_2_n_12, sub_352_2_n_13, sub_352_2_n_14, sub_352_2_n_15,
     sub_352_2_n_16, sub_352_2_n_20, sub_352_2_n_22, sub_352_2_n_23,
     sub_352_2_n_27, sub_352_2_n_28, sub_352_2_n_29, sub_352_2_n_30,
     sub_352_2_n_31, sub_352_2_n_32, sub_352_2_n_33, sub_352_2_n_36,
     sub_352_2_n_37, sub_352_2_n_38, sub_352_2_n_39, sub_352_2_n_40,
     sub_352_2_n_41, sub_352_2_n_42, sub_352_2_n_43, sub_352_2_n_44,
     sub_352_2_n_45, sub_352_2_n_46, sub_352_2_n_51, sub_352_2_n_52,
     sub_352_2_n_53, sub_352_2_n_54, sub_352_2_n_55, sub_352_2_n_57,
     sub_352_2_n_59, sub_352_2_n_60, sub_352_2_n_61, sub_352_2_n_63,
     sub_352_2_n_64, sub_352_2_n_65, sub_352_2_n_66, sub_352_2_n_70,
     sub_352_2_n_73, sub_352_2_n_74, sub_352_2_n_76, sub_352_2_n_77,
     sub_352_2_n_78, sub_352_2_n_81, sub_352_2_n_84, sub_352_2_n_86,
     sub_371_2_n_0, sub_371_2_n_1, sub_371_2_n_2, sub_371_2_n_3, sub_371_2_n_4,
     sub_371_2_n_5, sub_371_2_n_6, sub_371_2_n_7, sub_371_2_n_8, sub_371_2_n_9,
     sub_371_2_n_10, sub_371_2_n_11, sub_371_2_n_12, sub_371_2_n_13,
     sub_371_2_n_14, sub_371_2_n_15, sub_371_2_n_18, sub_371_2_n_19,
     sub_371_2_n_21, sub_371_2_n_23, sub_371_2_n_26, sub_371_2_n_27,
     sub_371_2_n_28, sub_371_2_n_29, sub_371_2_n_30, sub_371_2_n_31,
     sub_371_2_n_32, sub_371_2_n_33, sub_371_2_n_34, sub_371_2_n_35,
     sub_371_2_n_36, sub_371_2_n_38, sub_371_2_n_39, sub_371_2_n_40,
     sub_371_2_n_41, sub_371_2_n_42, sub_371_2_n_43, sub_371_2_n_44,
     sub_371_2_n_45, sub_371_2_n_46, sub_371_2_n_51, sub_371_2_n_52,
     sub_371_2_n_55, sub_371_2_n_56, sub_371_2_n_57, sub_371_2_n_58,
     sub_371_2_n_59, sub_371_2_n_60, sub_371_2_n_61, sub_371_2_n_62,
     sub_371_2_n_63, sub_371_2_n_64, sub_371_2_n_65, sub_371_2_n_67,
     sub_371_2_n_68, sub_371_2_n_69, sub_371_2_n_70, sub_371_2_n_71,
     sub_371_2_n_74, sub_371_2_n_75, sub_371_2_n_78, sub_371_2_n_79,
     sub_371_2_n_81, sub_371_2_n_82, sub_371_2_n_85, sub_371_2_n_88,
     sub_371_2_n_89, sub_371_2_n_92, sub_371_2_n_93, sub_371_2_n_96,
     sub_390_2_n_0, sub_390_2_n_1, sub_390_2_n_2, sub_390_2_n_3, sub_390_2_n_4,
     sub_390_2_n_5, sub_390_2_n_6, sub_390_2_n_7, sub_390_2_n_8, sub_390_2_n_9,
     sub_390_2_n_10, sub_390_2_n_11, sub_390_2_n_12, sub_390_2_n_13,
     sub_390_2_n_14, sub_390_2_n_17, sub_390_2_n_19, sub_390_2_n_21,
     sub_390_2_n_22, sub_390_2_n_23, sub_390_2_n_24, sub_390_2_n_25,
     sub_390_2_n_27, sub_390_2_n_28, sub_390_2_n_30, sub_390_2_n_31,
     sub_390_2_n_34, sub_390_2_n_35, sub_390_2_n_36, sub_390_2_n_37,
     sub_390_2_n_38, sub_390_2_n_41, sub_390_2_n_42, sub_390_2_n_43,
     sub_390_2_n_44, sub_390_2_n_45, sub_390_2_n_46, sub_390_2_n_47,
     sub_390_2_n_48, sub_390_2_n_49, sub_390_2_n_50, sub_390_2_n_52,
     sub_390_2_n_53, sub_390_2_n_54, sub_390_2_n_55, sub_390_2_n_56,
     sub_390_2_n_57, sub_390_2_n_58, sub_390_2_n_59, sub_390_2_n_63,
     sub_390_2_n_64, sub_390_2_n_65, sub_390_2_n_66, sub_390_2_n_67,
     sub_390_2_n_69, sub_390_2_n_70, sub_390_2_n_71, sub_390_2_n_73,
     sub_390_2_n_74, sub_390_2_n_76, sub_390_2_n_77, sub_390_2_n_79,
     sub_390_2_n_80, sub_390_2_n_81, sub_390_2_n_82, sub_390_2_n_83,
     sub_390_2_n_84, sub_390_2_n_85, sub_390_2_n_87, sub_390_2_n_88,
     sub_390_2_n_89, sub_390_2_n_91, sub_390_2_n_92, sub_390_2_n_95,
     sub_390_2_n_96, sub_390_2_n_98, sub_390_2_n_103, sub_390_2_n_107,
     sub_390_2_n_108, sub_409_2_n_0, sub_409_2_n_1, sub_409_2_n_2, sub_409_2_n_3,
     sub_409_2_n_4, sub_409_2_n_5, sub_409_2_n_7, sub_409_2_n_8, sub_409_2_n_9,
     sub_409_2_n_10, sub_409_2_n_11, sub_409_2_n_12, sub_409_2_n_15,
     sub_409_2_n_16, sub_409_2_n_17, sub_409_2_n_18, sub_409_2_n_22,
     sub_409_2_n_23, sub_409_2_n_24, sub_409_2_n_25, sub_409_2_n_26,
     sub_409_2_n_28, sub_409_2_n_29, sub_409_2_n_31, sub_409_2_n_34,
     sub_409_2_n_35, sub_409_2_n_37, sub_409_2_n_38, sub_409_2_n_39,
     sub_409_2_n_40, sub_409_2_n_41, sub_409_2_n_42, sub_409_2_n_43,
     sub_409_2_n_44, sub_409_2_n_45, sub_409_2_n_46, sub_409_2_n_47,
     sub_409_2_n_48, sub_409_2_n_49, sub_409_2_n_51, sub_409_2_n_52,
     sub_409_2_n_53, sub_409_2_n_54, sub_409_2_n_55, sub_409_2_n_56,
     sub_409_2_n_57, sub_409_2_n_59, sub_409_2_n_60, sub_409_2_n_61,
     sub_409_2_n_62, sub_409_2_n_63, sub_409_2_n_64, sub_409_2_n_65,
     sub_409_2_n_66, sub_409_2_n_67, sub_409_2_n_68, sub_409_2_n_69,
     sub_409_2_n_70, sub_409_2_n_71, sub_409_2_n_72, sub_409_2_n_73,
     sub_409_2_n_74, sub_409_2_n_75, sub_409_2_n_77, sub_409_2_n_78,
     sub_409_2_n_79, sub_409_2_n_80, sub_409_2_n_81, sub_409_2_n_83,
     sub_409_2_n_84, sub_409_2_n_85, sub_409_2_n_86, sub_409_2_n_88,
     sub_409_2_n_89, sub_409_2_n_90, sub_409_2_n_91, sub_409_2_n_97,
     sub_409_2_n_101, sub_409_2_n_102, sub_409_2_n_103, sub_428_2_n_0,
     sub_428_2_n_1, sub_428_2_n_2, sub_428_2_n_4, sub_428_2_n_5, sub_428_2_n_6,
     sub_428_2_n_7, sub_428_2_n_8, sub_428_2_n_9, sub_428_2_n_11, sub_428_2_n_12,
     sub_428_2_n_13, sub_428_2_n_14, sub_428_2_n_15, sub_428_2_n_17,
     sub_428_2_n_18, sub_428_2_n_19, sub_428_2_n_20, sub_428_2_n_21,
     sub_428_2_n_22, sub_428_2_n_26, sub_428_2_n_28, sub_428_2_n_29,
     sub_428_2_n_30, sub_428_2_n_31, sub_428_2_n_32, sub_428_2_n_33,
     sub_428_2_n_34, sub_428_2_n_36, sub_428_2_n_37, sub_428_2_n_38,
     sub_428_2_n_39, sub_428_2_n_40, sub_428_2_n_41, sub_428_2_n_43,
     sub_428_2_n_46, sub_428_2_n_47, sub_428_2_n_48, sub_428_2_n_49,
     sub_428_2_n_50, sub_428_2_n_51, sub_428_2_n_52, sub_428_2_n_54,
     sub_428_2_n_56, sub_428_2_n_57, sub_428_2_n_58, sub_428_2_n_59,
     sub_428_2_n_61, sub_428_2_n_62, sub_428_2_n_63, sub_428_2_n_64,
     sub_428_2_n_70, sub_428_2_n_71, sub_428_2_n_72, sub_428_2_n_74,
     sub_428_2_n_75, sub_428_2_n_76, sub_428_2_n_77, sub_428_2_n_78,
     sub_428_2_n_80, sub_428_2_n_81, sub_428_2_n_82, sub_428_2_n_83,
     sub_428_2_n_85, sub_428_2_n_87, sub_428_2_n_88, sub_428_2_n_89,
     sub_428_2_n_92, sub_428_2_n_93, sub_428_2_n_95, sub_428_2_n_99,
     sub_428_2_n_102, sub_428_2_n_103, sub_428_2_n_105, sub_428_2_n_109,
     sub_428_2_n_110, sub_428_2_n_111, sub_428_2_n_112, sub_428_2_n_113,
     sub_428_2_n_117, sub_428_2_n_118, sub_447_2_n_0, sub_447_2_n_1,
     sub_447_2_n_2, sub_447_2_n_3, sub_447_2_n_4, sub_447_2_n_5, sub_447_2_n_6,
     sub_447_2_n_7, sub_447_2_n_8, sub_447_2_n_9, sub_447_2_n_10, sub_447_2_n_11,
     sub_447_2_n_12, sub_447_2_n_13, sub_447_2_n_14, sub_447_2_n_15,
     sub_447_2_n_16, sub_447_2_n_17, sub_447_2_n_18, sub_447_2_n_19,
     sub_447_2_n_20, sub_447_2_n_23, sub_447_2_n_24, sub_447_2_n_25,
     sub_447_2_n_26, sub_447_2_n_27, sub_447_2_n_28, sub_447_2_n_29,
     sub_447_2_n_30, sub_447_2_n_34, sub_447_2_n_40, sub_447_2_n_41,
     sub_447_2_n_42, sub_447_2_n_43, sub_447_2_n_44, sub_447_2_n_45,
     sub_447_2_n_46, sub_447_2_n_47, sub_447_2_n_48, sub_447_2_n_49,
     sub_447_2_n_50, sub_447_2_n_55, sub_447_2_n_56, sub_447_2_n_57,
     sub_447_2_n_58, sub_447_2_n_59, sub_447_2_n_60, sub_447_2_n_61,
     sub_447_2_n_62, sub_447_2_n_64, sub_447_2_n_65, sub_447_2_n_66,
     sub_447_2_n_67, sub_447_2_n_68, sub_447_2_n_69, sub_447_2_n_74,
     sub_447_2_n_75, sub_447_2_n_76, sub_447_2_n_77, sub_447_2_n_78,
     sub_447_2_n_79, sub_447_2_n_80, sub_447_2_n_81, sub_447_2_n_82,
     sub_447_2_n_84, sub_447_2_n_85, sub_447_2_n_86, sub_447_2_n_87,
     sub_447_2_n_88, sub_447_2_n_89, sub_447_2_n_91, sub_447_2_n_92,
     sub_447_2_n_93, sub_447_2_n_94, sub_447_2_n_97, sub_447_2_n_99,
     sub_447_2_n_100, sub_447_2_n_105, sub_447_2_n_106, sub_447_2_n_107,
     sub_447_2_n_109, sub_447_2_n_111, sub_447_2_n_112, sub_447_2_n_114,
     sub_447_2_n_115, sub_447_2_n_116, sub_447_2_n_119, sub_447_2_n_120,
     sub_447_2_n_121, sub_447_2_n_123, sub_447_2_n_126, sub_447_2_n_127,
     sub_447_2_n_128, sub_447_2_n_132, sub_447_2_n_133, sub_447_2_n_134,
     sub_447_2_n_139, sub_466_2_n_0, sub_466_2_n_1, sub_466_2_n_2, sub_466_2_n_3,
     sub_466_2_n_4, sub_466_2_n_5, sub_466_2_n_6, sub_466_2_n_7, sub_466_2_n_8,
     sub_466_2_n_9, sub_466_2_n_10, sub_466_2_n_12, sub_466_2_n_13,
     sub_466_2_n_14, sub_466_2_n_15, sub_466_2_n_16, sub_466_2_n_17,
     sub_466_2_n_19, sub_466_2_n_24, sub_466_2_n_25, sub_466_2_n_26,
     sub_466_2_n_29, sub_466_2_n_31, sub_466_2_n_34, sub_466_2_n_35,
     sub_466_2_n_36, sub_466_2_n_39, sub_466_2_n_40, sub_466_2_n_41,
     sub_466_2_n_43, sub_466_2_n_44, sub_466_2_n_45, sub_466_2_n_46,
     sub_466_2_n_47, sub_466_2_n_48, sub_466_2_n_49, sub_466_2_n_50,
     sub_466_2_n_52, sub_466_2_n_53, sub_466_2_n_54, sub_466_2_n_55,
     sub_466_2_n_56, sub_466_2_n_57, sub_466_2_n_58, sub_466_2_n_60,
     sub_466_2_n_61, sub_466_2_n_62, sub_466_2_n_63, sub_466_2_n_64,
     sub_466_2_n_65, sub_466_2_n_66, sub_466_2_n_67, sub_466_2_n_68,
     sub_466_2_n_71, sub_466_2_n_73, sub_466_2_n_74, sub_466_2_n_75,
     sub_466_2_n_76, sub_466_2_n_77, sub_466_2_n_78, sub_466_2_n_79,
     sub_466_2_n_80, sub_466_2_n_81, sub_466_2_n_82, sub_466_2_n_83,
     sub_466_2_n_84, sub_466_2_n_85, sub_466_2_n_86, sub_466_2_n_87,
     sub_466_2_n_88, sub_466_2_n_89, sub_466_2_n_90, sub_466_2_n_91,
     sub_466_2_n_92, sub_466_2_n_93, sub_466_2_n_95, sub_466_2_n_96,
     sub_466_2_n_97, sub_466_2_n_98, sub_466_2_n_99, sub_466_2_n_100,
     sub_466_2_n_102, sub_466_2_n_103, sub_466_2_n_104, sub_466_2_n_105,
     sub_466_2_n_107, sub_466_2_n_110, sub_466_2_n_113, sub_466_2_n_117,
     sub_466_2_n_121, sub_466_2_n_122, sub_466_2_n_123, sub_466_2_n_127,
     sub_466_2_n_128, sub_466_2_n_129, sub_466_2_n_135, sub_485_2_n_0,
     sub_485_2_n_1, sub_485_2_n_2, sub_485_2_n_3, sub_485_2_n_4, sub_485_2_n_5,
     sub_485_2_n_6, sub_485_2_n_7, sub_485_2_n_8, sub_485_2_n_9, sub_485_2_n_10,
     sub_485_2_n_11, sub_485_2_n_12, sub_485_2_n_13, sub_485_2_n_14,
     sub_485_2_n_15, sub_485_2_n_16, sub_485_2_n_17, sub_485_2_n_18,
     sub_485_2_n_19, sub_485_2_n_20, sub_485_2_n_21, sub_485_2_n_22,
     sub_485_2_n_24, sub_485_2_n_27, sub_485_2_n_28, sub_485_2_n_30,
     sub_485_2_n_31, sub_485_2_n_32, sub_485_2_n_33, sub_485_2_n_34,
     sub_485_2_n_35, sub_485_2_n_36, sub_485_2_n_37, sub_485_2_n_38,
     sub_485_2_n_39, sub_485_2_n_40, sub_485_2_n_41, sub_485_2_n_42,
     sub_485_2_n_43, sub_485_2_n_45, sub_485_2_n_46, sub_485_2_n_47,
     sub_485_2_n_48, sub_485_2_n_49, sub_485_2_n_50, sub_485_2_n_51,
     sub_485_2_n_52, sub_485_2_n_54, sub_485_2_n_55, sub_485_2_n_56,
     sub_485_2_n_58, sub_485_2_n_60, sub_485_2_n_61, sub_485_2_n_62,
     sub_485_2_n_63, sub_485_2_n_66, sub_485_2_n_70, sub_485_2_n_71,
     sub_485_2_n_72, sub_485_2_n_73, sub_485_2_n_74, sub_485_2_n_75,
     sub_485_2_n_76, sub_485_2_n_77, sub_485_2_n_78, sub_485_2_n_79,
     sub_485_2_n_80, sub_485_2_n_82, sub_485_2_n_83, sub_485_2_n_84,
     sub_485_2_n_85, sub_485_2_n_86, sub_485_2_n_87, sub_485_2_n_88,
     sub_485_2_n_91, sub_485_2_n_92, sub_485_2_n_93, sub_485_2_n_94,
     sub_485_2_n_95, sub_485_2_n_97, sub_485_2_n_98, sub_485_2_n_100,
     sub_485_2_n_102, sub_485_2_n_103, sub_485_2_n_104, sub_485_2_n_108,
     sub_485_2_n_110, sub_485_2_n_115, sub_485_2_n_116, sub_485_2_n_117,
     sub_485_2_n_120, sub_485_2_n_121, sub_485_2_n_122, sub_485_2_n_126,
     sub_485_2_n_127, sub_485_2_n_128, sub_485_2_n_129, sub_485_2_n_133,
     sub_504_2_n_0, sub_504_2_n_1, sub_504_2_n_2, sub_504_2_n_3, sub_504_2_n_4,
     sub_504_2_n_5, sub_504_2_n_6, sub_504_2_n_7, sub_504_2_n_8, sub_504_2_n_9,
     sub_504_2_n_10, sub_504_2_n_11, sub_504_2_n_12, sub_504_2_n_13,
     sub_504_2_n_14, sub_504_2_n_15, sub_504_2_n_16, sub_504_2_n_17,
     sub_504_2_n_18, sub_504_2_n_19, sub_504_2_n_20, sub_504_2_n_22,
     sub_504_2_n_26, sub_504_2_n_28, sub_504_2_n_29, sub_504_2_n_30,
     sub_504_2_n_31, sub_504_2_n_32, sub_504_2_n_33, sub_504_2_n_34,
     sub_504_2_n_35, sub_504_2_n_36, sub_504_2_n_37, sub_504_2_n_38,
     sub_504_2_n_39, sub_504_2_n_40, sub_504_2_n_41, sub_504_2_n_42,
     sub_504_2_n_43, sub_504_2_n_44, sub_504_2_n_45, sub_504_2_n_46,
     sub_504_2_n_47, sub_504_2_n_48, sub_504_2_n_49, sub_504_2_n_50,
     sub_504_2_n_51, sub_504_2_n_52, sub_504_2_n_53, sub_504_2_n_54,
     sub_504_2_n_55, sub_504_2_n_56, sub_504_2_n_57, sub_504_2_n_58,
     sub_504_2_n_59, sub_504_2_n_60, sub_504_2_n_61, sub_504_2_n_62,
     sub_504_2_n_63, sub_504_2_n_64, sub_504_2_n_65, sub_504_2_n_67,
     sub_504_2_n_68, sub_504_2_n_69, sub_504_2_n_70, sub_504_2_n_71,
     sub_504_2_n_72, sub_504_2_n_73, sub_504_2_n_74, sub_504_2_n_75,
     sub_504_2_n_76, sub_504_2_n_77, sub_504_2_n_78, sub_504_2_n_81,
     sub_504_2_n_82, sub_504_2_n_83, sub_504_2_n_84, sub_504_2_n_86,
     sub_504_2_n_88, sub_504_2_n_89, sub_504_2_n_90, sub_504_2_n_91,
     sub_504_2_n_93, sub_504_2_n_95, sub_504_2_n_96, sub_504_2_n_97,
     sub_504_2_n_98, sub_504_2_n_99, sub_504_2_n_101, sub_504_2_n_102,
     sub_504_2_n_106, sub_504_2_n_107, sub_504_2_n_109, sub_504_2_n_115,
     sub_504_2_n_120, sub_504_2_n_121, sub_504_2_n_123, sub_504_2_n_127,
     sub_504_2_n_128, sub_504_2_n_129, sub_504_2_n_143, sub_504_2_n_147,
     sub_504_2_n_148, sub_523_2_n_0, sub_523_2_n_1, sub_523_2_n_2, sub_523_2_n_3,
     sub_523_2_n_4, sub_523_2_n_5, sub_523_2_n_6, sub_523_2_n_7, sub_523_2_n_8,
     sub_523_2_n_9, sub_523_2_n_10, sub_523_2_n_11, sub_523_2_n_12,
     sub_523_2_n_13, sub_523_2_n_14, sub_523_2_n_15, sub_523_2_n_16,
     sub_523_2_n_17, sub_523_2_n_18, sub_523_2_n_19, sub_523_2_n_20,
     sub_523_2_n_21, sub_523_2_n_22, sub_523_2_n_23, sub_523_2_n_24,
     sub_523_2_n_26, sub_523_2_n_27, sub_523_2_n_29, sub_523_2_n_31,
     sub_523_2_n_32, sub_523_2_n_33, sub_523_2_n_34, sub_523_2_n_35,
     sub_523_2_n_36, sub_523_2_n_37, sub_523_2_n_38, sub_523_2_n_39,
     sub_523_2_n_40, sub_523_2_n_41, sub_523_2_n_42, sub_523_2_n_43,
     sub_523_2_n_44, sub_523_2_n_45, sub_523_2_n_46, sub_523_2_n_47,
     sub_523_2_n_48, sub_523_2_n_49, sub_523_2_n_50, sub_523_2_n_52,
     sub_523_2_n_53, sub_523_2_n_54, sub_523_2_n_55, sub_523_2_n_56,
     sub_523_2_n_57, sub_523_2_n_58, sub_523_2_n_59, sub_523_2_n_60,
     sub_523_2_n_61, sub_523_2_n_62, sub_523_2_n_63, sub_523_2_n_64,
     sub_523_2_n_65, sub_523_2_n_67, sub_523_2_n_68, sub_523_2_n_69,
     sub_523_2_n_71, sub_523_2_n_74, sub_523_2_n_75, sub_523_2_n_76,
     sub_523_2_n_77, sub_523_2_n_78, sub_523_2_n_79, sub_523_2_n_80,
     sub_523_2_n_81, sub_523_2_n_82, sub_523_2_n_83, sub_523_2_n_84,
     sub_523_2_n_85, sub_523_2_n_86, sub_523_2_n_87, sub_523_2_n_88,
     sub_523_2_n_89, sub_523_2_n_90, sub_523_2_n_91, sub_523_2_n_92,
     sub_523_2_n_93, sub_523_2_n_94, sub_523_2_n_95, sub_523_2_n_96,
     sub_523_2_n_98, sub_523_2_n_100, sub_523_2_n_101, sub_523_2_n_102,
     sub_523_2_n_103, sub_523_2_n_105, sub_523_2_n_107, sub_523_2_n_111,
     sub_523_2_n_112, sub_523_2_n_118, sub_523_2_n_123, sub_523_2_n_124,
     sub_523_2_n_128, sub_523_2_n_129, sub_523_2_n_131, sub_523_2_n_136,
     sub_523_2_n_139, sub_542_2_n_0, sub_542_2_n_1, sub_542_2_n_2, sub_542_2_n_3,
     sub_542_2_n_4, sub_542_2_n_5, sub_542_2_n_6, sub_542_2_n_7, sub_542_2_n_8,
     sub_542_2_n_9, sub_542_2_n_10, sub_542_2_n_11, sub_542_2_n_12,
     sub_542_2_n_13, sub_542_2_n_14, sub_542_2_n_15, sub_542_2_n_16,
     sub_542_2_n_17, sub_542_2_n_18, sub_542_2_n_19, sub_542_2_n_21,
     sub_542_2_n_22, sub_542_2_n_23, sub_542_2_n_24, sub_542_2_n_25,
     sub_542_2_n_28, sub_542_2_n_31, sub_542_2_n_33, sub_542_2_n_34,
     sub_542_2_n_35, sub_542_2_n_36, sub_542_2_n_37, sub_542_2_n_38,
     sub_542_2_n_39, sub_542_2_n_40, sub_542_2_n_41, sub_542_2_n_42,
     sub_542_2_n_43, sub_542_2_n_44, sub_542_2_n_45, sub_542_2_n_46,
     sub_542_2_n_47, sub_542_2_n_48, sub_542_2_n_49, sub_542_2_n_50,
     sub_542_2_n_52, sub_542_2_n_53, sub_542_2_n_54, sub_542_2_n_55,
     sub_542_2_n_56, sub_542_2_n_57, sub_542_2_n_58, sub_542_2_n_59,
     sub_542_2_n_60, sub_542_2_n_61, sub_542_2_n_62, sub_542_2_n_63,
     sub_542_2_n_64, sub_542_2_n_65, sub_542_2_n_66, sub_542_2_n_67,
     sub_542_2_n_69, sub_542_2_n_71, sub_542_2_n_72, sub_542_2_n_73,
     sub_542_2_n_74, sub_542_2_n_75, sub_542_2_n_76, sub_542_2_n_77,
     sub_542_2_n_78, sub_542_2_n_79, sub_542_2_n_82, sub_542_2_n_83,
     sub_542_2_n_84, sub_542_2_n_85, sub_542_2_n_86, sub_542_2_n_87,
     sub_542_2_n_88, sub_542_2_n_89, sub_542_2_n_91, sub_542_2_n_92,
     sub_542_2_n_93, sub_542_2_n_94, sub_542_2_n_95, sub_542_2_n_96,
     sub_542_2_n_97, sub_542_2_n_99, sub_542_2_n_100, sub_542_2_n_101,
     sub_542_2_n_102, sub_542_2_n_103, sub_542_2_n_104, sub_542_2_n_107,
     sub_542_2_n_108, sub_542_2_n_109, sub_542_2_n_110, sub_542_2_n_111,
     sub_542_2_n_113, sub_542_2_n_116, sub_542_2_n_118, sub_542_2_n_125,
     sub_542_2_n_126, sub_542_2_n_128, sub_542_2_n_129, sub_542_2_n_132,
     sub_542_2_n_135, sub_542_2_n_137, sub_542_2_n_162, sub_561_2_n_0,
     sub_561_2_n_1, sub_561_2_n_2, sub_561_2_n_3, sub_561_2_n_4, sub_561_2_n_5,
     sub_561_2_n_6, sub_561_2_n_7, sub_561_2_n_8, sub_561_2_n_9, sub_561_2_n_10,
     sub_561_2_n_11, sub_561_2_n_12, sub_561_2_n_13, sub_561_2_n_14,
     sub_561_2_n_15, sub_561_2_n_16, sub_561_2_n_17, sub_561_2_n_18,
     sub_561_2_n_19, sub_561_2_n_20, sub_561_2_n_21, sub_561_2_n_22,
     sub_561_2_n_24, sub_561_2_n_25, sub_561_2_n_26, sub_561_2_n_27,
     sub_561_2_n_30, sub_561_2_n_31, sub_561_2_n_32, sub_561_2_n_33,
     sub_561_2_n_34, sub_561_2_n_36, sub_561_2_n_37, sub_561_2_n_38,
     sub_561_2_n_39, sub_561_2_n_40, sub_561_2_n_41, sub_561_2_n_42,
     sub_561_2_n_43, sub_561_2_n_44, sub_561_2_n_45, sub_561_2_n_46,
     sub_561_2_n_47, sub_561_2_n_48, sub_561_2_n_49, sub_561_2_n_50,
     sub_561_2_n_51, sub_561_2_n_52, sub_561_2_n_55, sub_561_2_n_56,
     sub_561_2_n_57, sub_561_2_n_58, sub_561_2_n_59, sub_561_2_n_60,
     sub_561_2_n_61, sub_561_2_n_62, sub_561_2_n_63, sub_561_2_n_64,
     sub_561_2_n_65, sub_561_2_n_66, sub_561_2_n_67, sub_561_2_n_68,
     sub_561_2_n_70, sub_561_2_n_71, sub_561_2_n_72, sub_561_2_n_73,
     sub_561_2_n_74, sub_561_2_n_75, sub_561_2_n_76, sub_561_2_n_77,
     sub_561_2_n_78, sub_561_2_n_80, sub_561_2_n_83, sub_561_2_n_85,
     sub_561_2_n_86, sub_561_2_n_87, sub_561_2_n_88, sub_561_2_n_89,
     sub_561_2_n_90, sub_561_2_n_91, sub_561_2_n_92, sub_561_2_n_95,
     sub_561_2_n_96, sub_561_2_n_97, sub_561_2_n_98, sub_561_2_n_99,
     sub_561_2_n_100, sub_561_2_n_101, sub_561_2_n_102, sub_561_2_n_104,
     sub_561_2_n_105, sub_561_2_n_106, sub_561_2_n_107, sub_561_2_n_109,
     sub_561_2_n_110, sub_561_2_n_111, sub_561_2_n_112, sub_561_2_n_113,
     sub_561_2_n_115, sub_561_2_n_117, sub_561_2_n_119, sub_561_2_n_121,
     sub_561_2_n_122, sub_561_2_n_132, sub_561_2_n_133, sub_561_2_n_137,
     sub_561_2_n_138, sub_561_2_n_139, sub_561_2_n_143, sub_561_2_n_145,
     sub_561_2_n_152, sub_561_2_n_153, sub_561_2_n_163, sub_561_2_n_172,
     sub_580_2_n_0, sub_580_2_n_1, sub_580_2_n_2, sub_580_2_n_3, sub_580_2_n_4,
     sub_580_2_n_5, sub_580_2_n_6, sub_580_2_n_7, sub_580_2_n_8, sub_580_2_n_9,
     sub_580_2_n_10, sub_580_2_n_11, sub_580_2_n_12, sub_580_2_n_13,
     sub_580_2_n_14, sub_580_2_n_15, sub_580_2_n_16, sub_580_2_n_17,
     sub_580_2_n_18, sub_580_2_n_19, sub_580_2_n_20, sub_580_2_n_21,
     sub_580_2_n_22, sub_580_2_n_23, sub_580_2_n_24, sub_580_2_n_25,
     sub_580_2_n_26, sub_580_2_n_27, sub_580_2_n_28, sub_580_2_n_29,
     sub_580_2_n_30, sub_580_2_n_31, sub_580_2_n_32, sub_580_2_n_33,
     sub_580_2_n_37, sub_580_2_n_40, sub_580_2_n_41, sub_580_2_n_42,
     sub_580_2_n_43, sub_580_2_n_44, sub_580_2_n_45, sub_580_2_n_46,
     sub_580_2_n_47, sub_580_2_n_48, sub_580_2_n_49, sub_580_2_n_50,
     sub_580_2_n_51, sub_580_2_n_52, sub_580_2_n_53, sub_580_2_n_54,
     sub_580_2_n_55, sub_580_2_n_56, sub_580_2_n_57, sub_580_2_n_59,
     sub_580_2_n_60, sub_580_2_n_61, sub_580_2_n_62, sub_580_2_n_63,
     sub_580_2_n_64, sub_580_2_n_65, sub_580_2_n_66, sub_580_2_n_67,
     sub_580_2_n_68, sub_580_2_n_69, sub_580_2_n_70, sub_580_2_n_71,
     sub_580_2_n_72, sub_580_2_n_73, sub_580_2_n_74, sub_580_2_n_75,
     sub_580_2_n_76, sub_580_2_n_77, sub_580_2_n_78, sub_580_2_n_79,
     sub_580_2_n_80, sub_580_2_n_81, sub_580_2_n_82, sub_580_2_n_83,
     sub_580_2_n_85, sub_580_2_n_87, sub_580_2_n_88, sub_580_2_n_89,
     sub_580_2_n_90, sub_580_2_n_91, sub_580_2_n_92, sub_580_2_n_93,
     sub_580_2_n_94, sub_580_2_n_95, sub_580_2_n_96, sub_580_2_n_97,
     sub_580_2_n_98, sub_580_2_n_99, sub_580_2_n_100, sub_580_2_n_101,
     sub_580_2_n_102, sub_580_2_n_103, sub_580_2_n_104, sub_580_2_n_105,
     sub_580_2_n_106, sub_580_2_n_107, sub_580_2_n_108, sub_580_2_n_109,
     sub_580_2_n_110, sub_580_2_n_111, sub_580_2_n_113, sub_580_2_n_114,
     sub_580_2_n_115, sub_580_2_n_117, sub_580_2_n_118, sub_580_2_n_121,
     sub_580_2_n_123, sub_580_2_n_125, sub_580_2_n_127, sub_580_2_n_128,
     sub_580_2_n_130, sub_580_2_n_131, sub_580_2_n_133, sub_580_2_n_137,
     sub_580_2_n_138, sub_580_2_n_139, sub_580_2_n_140, sub_580_2_n_145,
     sub_580_2_n_149, sub_580_2_n_153, sub_580_2_n_154, sub_580_2_n_160,
     sub_580_2_n_170, sub_580_2_n_174, sub_599_2_n_0, sub_599_2_n_1,
     sub_599_2_n_2, sub_599_2_n_3, sub_599_2_n_4, sub_599_2_n_5, sub_599_2_n_6,
     sub_599_2_n_7, sub_599_2_n_8, sub_599_2_n_9, sub_599_2_n_10, sub_599_2_n_11,
     sub_599_2_n_12, sub_599_2_n_13, sub_599_2_n_14, sub_599_2_n_15,
     sub_599_2_n_16, sub_599_2_n_17, sub_599_2_n_18, sub_599_2_n_19,
     sub_599_2_n_20, sub_599_2_n_21, sub_599_2_n_22, sub_599_2_n_23,
     sub_599_2_n_24, sub_599_2_n_26, sub_599_2_n_27, sub_599_2_n_28,
     sub_599_2_n_29, sub_599_2_n_30, sub_599_2_n_31, sub_599_2_n_32,
     sub_599_2_n_33, sub_599_2_n_34, sub_599_2_n_35, sub_599_2_n_36,
     sub_599_2_n_37, sub_599_2_n_38, sub_599_2_n_39, sub_599_2_n_40,
     sub_599_2_n_41, sub_599_2_n_43, sub_599_2_n_44, sub_599_2_n_45,
     sub_599_2_n_46, sub_599_2_n_48, sub_599_2_n_49, sub_599_2_n_50,
     sub_599_2_n_51, sub_599_2_n_52, sub_599_2_n_53, sub_599_2_n_54,
     sub_599_2_n_55, sub_599_2_n_56, sub_599_2_n_57, sub_599_2_n_58,
     sub_599_2_n_59, sub_599_2_n_60, sub_599_2_n_61, sub_599_2_n_62,
     sub_599_2_n_63, sub_599_2_n_64, sub_599_2_n_65, sub_599_2_n_68,
     sub_599_2_n_69, sub_599_2_n_70, sub_599_2_n_71, sub_599_2_n_72,
     sub_599_2_n_73, sub_599_2_n_74, sub_599_2_n_75, sub_599_2_n_76,
     sub_599_2_n_77, sub_599_2_n_78, sub_599_2_n_79, sub_599_2_n_80,
     sub_599_2_n_81, sub_599_2_n_83, sub_599_2_n_84, sub_599_2_n_85,
     sub_599_2_n_86, sub_599_2_n_87, sub_599_2_n_90, sub_599_2_n_91,
     sub_599_2_n_92, sub_599_2_n_93, sub_599_2_n_94, sub_599_2_n_95,
     sub_599_2_n_96, sub_599_2_n_97, sub_599_2_n_98, sub_599_2_n_99,
     sub_599_2_n_100, sub_599_2_n_101, sub_599_2_n_104, sub_599_2_n_105,
     sub_599_2_n_106, sub_599_2_n_107, sub_599_2_n_108, sub_599_2_n_109,
     sub_599_2_n_110, sub_599_2_n_111, sub_599_2_n_112, sub_599_2_n_113,
     sub_599_2_n_114, sub_599_2_n_115, sub_599_2_n_116, sub_599_2_n_117,
     sub_599_2_n_118, sub_599_2_n_119, sub_599_2_n_120, sub_599_2_n_121,
     sub_599_2_n_122, sub_599_2_n_123, sub_599_2_n_125, sub_599_2_n_127,
     sub_599_2_n_129, sub_599_2_n_130, sub_599_2_n_131, sub_599_2_n_132,
     sub_599_2_n_134, sub_599_2_n_135, sub_599_2_n_136, sub_599_2_n_139,
     sub_599_2_n_140, sub_599_2_n_141, sub_599_2_n_145, sub_599_2_n_149,
     sub_599_2_n_151, sub_599_2_n_152, sub_599_2_n_153, sub_599_2_n_158,
     sub_599_2_n_159, sub_599_2_n_160, sub_599_2_n_161, sub_599_2_n_168,
     sub_599_2_n_169, sub_599_2_n_170, sub_599_2_n_171, sub_618_2_n_0,
     sub_618_2_n_1, sub_618_2_n_2, sub_618_2_n_3, sub_618_2_n_4, sub_618_2_n_5,
     sub_618_2_n_6, sub_618_2_n_7, sub_618_2_n_8, sub_618_2_n_9, sub_618_2_n_10,
     sub_618_2_n_11, sub_618_2_n_12, sub_618_2_n_13, sub_618_2_n_14,
     sub_618_2_n_15, sub_618_2_n_16, sub_618_2_n_17, sub_618_2_n_18,
     sub_618_2_n_19, sub_618_2_n_20, sub_618_2_n_22, sub_618_2_n_23,
     sub_618_2_n_24, sub_618_2_n_25, sub_618_2_n_26, sub_618_2_n_27,
     sub_618_2_n_28, sub_618_2_n_29, sub_618_2_n_30, sub_618_2_n_31,
     sub_618_2_n_32, sub_618_2_n_33, sub_618_2_n_42, sub_618_2_n_43,
     sub_618_2_n_44, sub_618_2_n_45, sub_618_2_n_46, sub_618_2_n_47,
     sub_618_2_n_48, sub_618_2_n_49, sub_618_2_n_50, sub_618_2_n_51,
     sub_618_2_n_52, sub_618_2_n_53, sub_618_2_n_54, sub_618_2_n_55,
     sub_618_2_n_56, sub_618_2_n_57, sub_618_2_n_58, sub_618_2_n_59,
     sub_618_2_n_60, sub_618_2_n_61, sub_618_2_n_62, sub_618_2_n_63,
     sub_618_2_n_64, sub_618_2_n_65, sub_618_2_n_66, sub_618_2_n_67,
     sub_618_2_n_68, sub_618_2_n_69, sub_618_2_n_70, sub_618_2_n_71,
     sub_618_2_n_72, sub_618_2_n_73, sub_618_2_n_74, sub_618_2_n_75,
     sub_618_2_n_76, sub_618_2_n_77, sub_618_2_n_78, sub_618_2_n_79,
     sub_618_2_n_80, sub_618_2_n_81, sub_618_2_n_82, sub_618_2_n_83,
     sub_618_2_n_84, sub_618_2_n_86, sub_618_2_n_87, sub_618_2_n_88,
     sub_618_2_n_89, sub_618_2_n_90, sub_618_2_n_91, sub_618_2_n_92,
     sub_618_2_n_93, sub_618_2_n_94, sub_618_2_n_95, sub_618_2_n_97,
     sub_618_2_n_99, sub_618_2_n_100, sub_618_2_n_101, sub_618_2_n_102,
     sub_618_2_n_103, sub_618_2_n_104, sub_618_2_n_107, sub_618_2_n_108,
     sub_618_2_n_109, sub_618_2_n_110, sub_618_2_n_111, sub_618_2_n_112,
     sub_618_2_n_113, sub_618_2_n_114, sub_618_2_n_115, sub_618_2_n_116,
     sub_618_2_n_117, sub_618_2_n_118, sub_618_2_n_120, sub_618_2_n_121,
     sub_618_2_n_122, sub_618_2_n_123, sub_618_2_n_124, sub_618_2_n_126,
     sub_618_2_n_127, sub_618_2_n_129, sub_618_2_n_130, sub_618_2_n_131,
     sub_618_2_n_132, sub_618_2_n_134, sub_618_2_n_136, sub_618_2_n_137,
     sub_618_2_n_138, sub_618_2_n_139, sub_618_2_n_141, sub_618_2_n_142,
     sub_618_2_n_146, sub_618_2_n_152, sub_618_2_n_160, sub_618_2_n_161,
     sub_618_2_n_170, sub_618_2_n_174, sub_618_2_n_175, sub_618_2_n_181,
     sub_637_2_n_0, sub_637_2_n_1, sub_637_2_n_2, sub_637_2_n_3, sub_637_2_n_4,
     sub_637_2_n_5, sub_637_2_n_6, sub_637_2_n_7, sub_637_2_n_8, sub_637_2_n_9,
     sub_637_2_n_10, sub_637_2_n_11, sub_637_2_n_12, sub_637_2_n_13,
     sub_637_2_n_14, sub_637_2_n_15, sub_637_2_n_16, sub_637_2_n_17,
     sub_637_2_n_18, sub_637_2_n_19, sub_637_2_n_20, sub_637_2_n_21,
     sub_637_2_n_22, sub_637_2_n_23, sub_637_2_n_25, sub_637_2_n_28,
     sub_637_2_n_29, sub_637_2_n_30, sub_637_2_n_32, sub_637_2_n_33,
     sub_637_2_n_34, sub_637_2_n_35, sub_637_2_n_36, sub_637_2_n_37,
     sub_637_2_n_38, sub_637_2_n_39, sub_637_2_n_40, sub_637_2_n_41,
     sub_637_2_n_42, sub_637_2_n_43, sub_637_2_n_44, sub_637_2_n_45,
     sub_637_2_n_46, sub_637_2_n_47, sub_637_2_n_48, sub_637_2_n_49,
     sub_637_2_n_50, sub_637_2_n_51, sub_637_2_n_52, sub_637_2_n_53,
     sub_637_2_n_54, sub_637_2_n_55, sub_637_2_n_56, sub_637_2_n_57,
     sub_637_2_n_58, sub_637_2_n_59, sub_637_2_n_60, sub_637_2_n_61,
     sub_637_2_n_62, sub_637_2_n_63, sub_637_2_n_64, sub_637_2_n_65,
     sub_637_2_n_66, sub_637_2_n_67, sub_637_2_n_68, sub_637_2_n_69,
     sub_637_2_n_70, sub_637_2_n_71, sub_637_2_n_72, sub_637_2_n_73,
     sub_637_2_n_74, sub_637_2_n_75, sub_637_2_n_76, sub_637_2_n_78,
     sub_637_2_n_79, sub_637_2_n_80, sub_637_2_n_81, sub_637_2_n_82,
     sub_637_2_n_83, sub_637_2_n_84, sub_637_2_n_85, sub_637_2_n_86,
     sub_637_2_n_87, sub_637_2_n_88, sub_637_2_n_92, sub_637_2_n_93,
     sub_637_2_n_94, sub_637_2_n_95, sub_637_2_n_96, sub_637_2_n_97,
     sub_637_2_n_98, sub_637_2_n_99, sub_637_2_n_100, sub_637_2_n_101,
     sub_637_2_n_102, sub_637_2_n_103, sub_637_2_n_104, sub_637_2_n_105,
     sub_637_2_n_106, sub_637_2_n_109, sub_637_2_n_110, sub_637_2_n_111,
     sub_637_2_n_112, sub_637_2_n_113, sub_637_2_n_114, sub_637_2_n_115,
     sub_637_2_n_116, sub_637_2_n_117, sub_637_2_n_118, sub_637_2_n_119,
     sub_637_2_n_121, sub_637_2_n_122, sub_637_2_n_123, sub_637_2_n_124,
     sub_637_2_n_125, sub_637_2_n_126, sub_637_2_n_128, sub_637_2_n_132,
     sub_637_2_n_134, sub_637_2_n_135, sub_637_2_n_136, sub_637_2_n_137,
     sub_637_2_n_138, sub_637_2_n_140, sub_637_2_n_141, sub_637_2_n_143,
     sub_637_2_n_144, sub_637_2_n_145, sub_637_2_n_146, sub_637_2_n_148,
     sub_637_2_n_149, sub_637_2_n_150, sub_637_2_n_153, sub_637_2_n_157,
     sub_637_2_n_158, sub_637_2_n_162, sub_637_2_n_163, sub_637_2_n_164,
     sub_637_2_n_168, sub_637_2_n_169, sub_637_2_n_173, sub_637_2_n_174,
     sub_637_2_n_175, sub_637_2_n_176, sub_637_2_n_180, sub_637_2_n_188,
     sub_637_2_n_189, sub_656_2_n_0, sub_656_2_n_1, sub_656_2_n_2, sub_656_2_n_3,
     sub_656_2_n_4, sub_656_2_n_5, sub_656_2_n_6, sub_656_2_n_7, sub_656_2_n_8,
     sub_656_2_n_9, sub_656_2_n_10, sub_656_2_n_11, sub_656_2_n_12,
     sub_656_2_n_13, sub_656_2_n_14, sub_656_2_n_15, sub_656_2_n_16,
     sub_656_2_n_17, sub_656_2_n_18, sub_656_2_n_19, sub_656_2_n_20,
     sub_656_2_n_23, sub_656_2_n_24, sub_656_2_n_25, sub_656_2_n_26,
     sub_656_2_n_27, sub_656_2_n_29, sub_656_2_n_32, sub_656_2_n_33,
     sub_656_2_n_34, sub_656_2_n_35, sub_656_2_n_37, sub_656_2_n_38,
     sub_656_2_n_39, sub_656_2_n_40, sub_656_2_n_41, sub_656_2_n_42,
     sub_656_2_n_43, sub_656_2_n_44, sub_656_2_n_45, sub_656_2_n_46,
     sub_656_2_n_47, sub_656_2_n_48, sub_656_2_n_49, sub_656_2_n_50,
     sub_656_2_n_51, sub_656_2_n_52, sub_656_2_n_53, sub_656_2_n_54,
     sub_656_2_n_55, sub_656_2_n_56, sub_656_2_n_57, sub_656_2_n_58,
     sub_656_2_n_59, sub_656_2_n_60, sub_656_2_n_61, sub_656_2_n_62,
     sub_656_2_n_63, sub_656_2_n_64, sub_656_2_n_65, sub_656_2_n_66,
     sub_656_2_n_67, sub_656_2_n_68, sub_656_2_n_69, sub_656_2_n_70,
     sub_656_2_n_71, sub_656_2_n_72, sub_656_2_n_73, sub_656_2_n_74,
     sub_656_2_n_75, sub_656_2_n_76, sub_656_2_n_77, sub_656_2_n_78,
     sub_656_2_n_79, sub_656_2_n_80, sub_656_2_n_81, sub_656_2_n_82,
     sub_656_2_n_83, sub_656_2_n_84, sub_656_2_n_85, sub_656_2_n_86,
     sub_656_2_n_87, sub_656_2_n_88, sub_656_2_n_89, sub_656_2_n_90,
     sub_656_2_n_91, sub_656_2_n_92, sub_656_2_n_93, sub_656_2_n_94,
     sub_656_2_n_95, sub_656_2_n_98, sub_656_2_n_99, sub_656_2_n_100,
     sub_656_2_n_101, sub_656_2_n_102, sub_656_2_n_103, sub_656_2_n_104,
     sub_656_2_n_105, sub_656_2_n_106, sub_656_2_n_107, sub_656_2_n_108,
     sub_656_2_n_109, sub_656_2_n_110, sub_656_2_n_111, sub_656_2_n_112,
     sub_656_2_n_113, sub_656_2_n_114, sub_656_2_n_115, sub_656_2_n_116,
     sub_656_2_n_117, sub_656_2_n_118, sub_656_2_n_119, sub_656_2_n_120,
     sub_656_2_n_121, sub_656_2_n_122, sub_656_2_n_123, sub_656_2_n_124,
     sub_656_2_n_125, sub_656_2_n_126, sub_656_2_n_127, sub_656_2_n_128,
     sub_656_2_n_129, sub_656_2_n_130, sub_656_2_n_132, sub_656_2_n_133,
     sub_656_2_n_134, sub_656_2_n_135, sub_656_2_n_136, sub_656_2_n_138,
     sub_656_2_n_139, sub_656_2_n_142, sub_656_2_n_143, sub_656_2_n_144,
     sub_656_2_n_145, sub_656_2_n_147, sub_656_2_n_148, sub_656_2_n_151,
     sub_656_2_n_152, sub_656_2_n_157, sub_656_2_n_159, sub_656_2_n_164,
     sub_656_2_n_165, sub_656_2_n_168, sub_656_2_n_173, sub_656_2_n_174,
     sub_656_2_n_183, sub_656_2_n_187, sub_656_2_n_188, sub_675_2_n_0,
     sub_675_2_n_1, sub_675_2_n_2, sub_675_2_n_3, sub_675_2_n_4, sub_675_2_n_5,
     sub_675_2_n_6, sub_675_2_n_7, sub_675_2_n_8, sub_675_2_n_9, sub_675_2_n_10,
     sub_675_2_n_11, sub_675_2_n_12, sub_675_2_n_13, sub_675_2_n_14,
     sub_675_2_n_15, sub_675_2_n_16, sub_675_2_n_17, sub_675_2_n_19,
     sub_675_2_n_21, sub_675_2_n_22, sub_675_2_n_24, sub_675_2_n_25,
     sub_675_2_n_26, sub_675_2_n_28, sub_675_2_n_29, sub_675_2_n_30,
     sub_675_2_n_31, sub_675_2_n_32, sub_675_2_n_33, sub_675_2_n_34,
     sub_675_2_n_35, sub_675_2_n_36, sub_675_2_n_37, sub_675_2_n_38,
     sub_675_2_n_39, sub_675_2_n_40, sub_675_2_n_41, sub_675_2_n_42,
     sub_675_2_n_43, sub_675_2_n_44, sub_675_2_n_45, sub_675_2_n_46,
     sub_675_2_n_47, sub_675_2_n_48, sub_675_2_n_49, sub_675_2_n_50,
     sub_675_2_n_51, sub_675_2_n_52, sub_675_2_n_53, sub_675_2_n_54,
     sub_675_2_n_55, sub_675_2_n_56, sub_675_2_n_57, sub_675_2_n_58,
     sub_675_2_n_59, sub_675_2_n_60, sub_675_2_n_61, sub_675_2_n_62,
     sub_675_2_n_63, sub_675_2_n_64, sub_675_2_n_65, sub_675_2_n_66,
     sub_675_2_n_67, sub_675_2_n_68, sub_675_2_n_69, sub_675_2_n_70,
     sub_675_2_n_72, sub_675_2_n_73, sub_675_2_n_74, sub_675_2_n_75,
     sub_675_2_n_76, sub_675_2_n_77, sub_675_2_n_78, sub_675_2_n_79,
     sub_675_2_n_80, sub_675_2_n_81, sub_675_2_n_82, sub_675_2_n_83,
     sub_675_2_n_84, sub_675_2_n_85, sub_675_2_n_87, sub_675_2_n_89,
     sub_675_2_n_90, sub_675_2_n_91, sub_675_2_n_92, sub_675_2_n_93,
     sub_675_2_n_94, sub_675_2_n_95, sub_675_2_n_96, sub_675_2_n_97,
     sub_675_2_n_98, sub_675_2_n_99, sub_675_2_n_100, sub_675_2_n_101,
     sub_675_2_n_102, sub_675_2_n_103, sub_675_2_n_104, sub_675_2_n_105,
     sub_675_2_n_106, sub_675_2_n_107, sub_675_2_n_108, sub_675_2_n_109,
     sub_675_2_n_110, sub_675_2_n_111, sub_675_2_n_115, sub_675_2_n_116,
     sub_675_2_n_117, sub_675_2_n_118, sub_675_2_n_119, sub_675_2_n_121,
     sub_675_2_n_123, sub_675_2_n_125, sub_675_2_n_126, sub_675_2_n_127,
     sub_675_2_n_128, sub_675_2_n_129, sub_675_2_n_130, sub_675_2_n_131,
     sub_675_2_n_132, sub_675_2_n_133, sub_675_2_n_134, sub_675_2_n_135,
     sub_675_2_n_137, sub_675_2_n_138, sub_675_2_n_139, sub_675_2_n_140,
     sub_675_2_n_141, sub_675_2_n_143, sub_675_2_n_144, sub_675_2_n_146,
     sub_675_2_n_147, sub_675_2_n_148, sub_675_2_n_149, sub_675_2_n_151,
     sub_675_2_n_152, sub_675_2_n_154, sub_675_2_n_155, sub_675_2_n_156,
     sub_675_2_n_159, sub_675_2_n_165, sub_675_2_n_166, sub_675_2_n_168,
     sub_675_2_n_169, sub_675_2_n_170, sub_675_2_n_174, sub_675_2_n_175,
     sub_675_2_n_176, sub_675_2_n_181, sub_675_2_n_184, sub_675_2_n_188,
     sub_675_2_n_189, sub_675_2_n_196, sub_675_2_n_197, sub_675_2_n_198,
     sub_675_2_n_199, sub_675_2_n_207, sub_694_2_n_0, sub_694_2_n_1,
     sub_694_2_n_2, sub_694_2_n_3, sub_694_2_n_4, sub_694_2_n_5, sub_694_2_n_6,
     sub_694_2_n_7, sub_694_2_n_9, sub_694_2_n_10, sub_694_2_n_11,
     sub_694_2_n_12, sub_694_2_n_13, sub_694_2_n_14, sub_694_2_n_15,
     sub_694_2_n_16, sub_694_2_n_17, sub_694_2_n_18, sub_694_2_n_19,
     sub_694_2_n_20, sub_694_2_n_21, sub_694_2_n_22, sub_694_2_n_23,
     sub_694_2_n_24, sub_694_2_n_25, sub_694_2_n_26, sub_694_2_n_27,
     sub_694_2_n_28, sub_694_2_n_29, sub_694_2_n_30, sub_694_2_n_31,
     sub_694_2_n_32, sub_694_2_n_33, sub_694_2_n_34, sub_694_2_n_35,
     sub_694_2_n_36, sub_694_2_n_37, sub_694_2_n_38, sub_694_2_n_39,
     sub_694_2_n_40, sub_694_2_n_41, sub_694_2_n_42, sub_694_2_n_43,
     sub_694_2_n_44, sub_694_2_n_45, sub_694_2_n_46, sub_694_2_n_47,
     sub_694_2_n_48, sub_694_2_n_49, sub_694_2_n_50, sub_694_2_n_51,
     sub_694_2_n_52, sub_694_2_n_53, sub_694_2_n_54, sub_694_2_n_55,
     sub_694_2_n_56, sub_694_2_n_57, sub_694_2_n_58, sub_694_2_n_59,
     sub_694_2_n_60, sub_694_2_n_61, sub_694_2_n_62, sub_694_2_n_63,
     sub_694_2_n_64, sub_694_2_n_65, sub_694_2_n_66, sub_694_2_n_67,
     sub_694_2_n_68, sub_694_2_n_69, sub_694_2_n_70, sub_694_2_n_71,
     sub_694_2_n_72, sub_694_2_n_73, sub_694_2_n_74, sub_694_2_n_75,
     sub_694_2_n_76, sub_694_2_n_78, sub_694_2_n_79, sub_694_2_n_80,
     sub_694_2_n_81, sub_694_2_n_82, sub_694_2_n_83, sub_694_2_n_84,
     sub_694_2_n_85, sub_694_2_n_86, sub_694_2_n_87, sub_694_2_n_88,
     sub_694_2_n_89, sub_694_2_n_90, sub_694_2_n_91, sub_694_2_n_92,
     sub_694_2_n_93, sub_694_2_n_94, sub_694_2_n_95, sub_694_2_n_96,
     sub_694_2_n_97, sub_694_2_n_98, sub_694_2_n_99, sub_694_2_n_100,
     sub_694_2_n_102, sub_694_2_n_103, sub_694_2_n_104, sub_694_2_n_105,
     sub_694_2_n_106, sub_694_2_n_107, sub_694_2_n_108, sub_694_2_n_109,
     sub_694_2_n_110, sub_694_2_n_111, sub_694_2_n_112, sub_694_2_n_113,
     sub_694_2_n_114, sub_694_2_n_115, sub_694_2_n_116, sub_694_2_n_117,
     sub_694_2_n_118, sub_694_2_n_119, sub_694_2_n_120, sub_694_2_n_121,
     sub_694_2_n_122, sub_694_2_n_123, sub_694_2_n_124, sub_694_2_n_126,
     sub_694_2_n_127, sub_694_2_n_128, sub_694_2_n_129, sub_694_2_n_130,
     sub_694_2_n_132, sub_694_2_n_133, sub_694_2_n_135, sub_694_2_n_136,
     sub_694_2_n_137, sub_694_2_n_138, sub_694_2_n_142, sub_694_2_n_143,
     sub_694_2_n_145, sub_694_2_n_146, sub_694_2_n_147, sub_694_2_n_150,
     sub_694_2_n_151, sub_694_2_n_152, sub_694_2_n_155, sub_694_2_n_156,
     sub_694_2_n_157, sub_694_2_n_158, sub_694_2_n_159, sub_694_2_n_160,
     sub_694_2_n_164, sub_694_2_n_165, sub_694_2_n_166, sub_694_2_n_168,
     sub_694_2_n_169, sub_694_2_n_170, sub_694_2_n_171, sub_694_2_n_175,
     sub_694_2_n_176, sub_694_2_n_182, sub_694_2_n_183, sub_694_2_n_184,
     sub_694_2_n_187, sub_694_2_n_188, sub_694_2_n_192, sub_694_2_n_196,
     sub_713_2_n_0, sub_713_2_n_1, sub_713_2_n_2, sub_713_2_n_4, sub_713_2_n_5,
     sub_713_2_n_6, sub_713_2_n_7, sub_713_2_n_8, sub_713_2_n_9, sub_713_2_n_10,
     sub_713_2_n_11, sub_713_2_n_12, sub_713_2_n_13, sub_713_2_n_14,
     sub_713_2_n_15, sub_713_2_n_16, sub_713_2_n_17, sub_713_2_n_18,
     sub_713_2_n_19, sub_713_2_n_20, sub_713_2_n_21, sub_713_2_n_22,
     sub_713_2_n_23, sub_713_2_n_24, sub_713_2_n_25, sub_713_2_n_26,
     sub_713_2_n_27, sub_713_2_n_28, sub_713_2_n_29, sub_713_2_n_30,
     sub_713_2_n_31, sub_713_2_n_32, sub_713_2_n_33, sub_713_2_n_34,
     sub_713_2_n_35, sub_713_2_n_36, sub_713_2_n_37, sub_713_2_n_38,
     sub_713_2_n_39, sub_713_2_n_40, sub_713_2_n_41, sub_713_2_n_42,
     sub_713_2_n_43, sub_713_2_n_44, sub_713_2_n_45, sub_713_2_n_46,
     sub_713_2_n_47, sub_713_2_n_48, sub_713_2_n_49, sub_713_2_n_50,
     sub_713_2_n_51, sub_713_2_n_52, sub_713_2_n_53, sub_713_2_n_54,
     sub_713_2_n_55, sub_713_2_n_56, sub_713_2_n_57, sub_713_2_n_58,
     sub_713_2_n_59, sub_713_2_n_60, sub_713_2_n_61, sub_713_2_n_62,
     sub_713_2_n_63, sub_713_2_n_64, sub_713_2_n_65, sub_713_2_n_66,
     sub_713_2_n_67, sub_713_2_n_68, sub_713_2_n_69, sub_713_2_n_70,
     sub_713_2_n_71, sub_713_2_n_72, sub_713_2_n_73, sub_713_2_n_74,
     sub_713_2_n_75, sub_713_2_n_76, sub_713_2_n_77, sub_713_2_n_78,
     sub_713_2_n_80, sub_713_2_n_81, sub_713_2_n_82, sub_713_2_n_83,
     sub_713_2_n_84, sub_713_2_n_85, sub_713_2_n_86, sub_713_2_n_87,
     sub_713_2_n_88, sub_713_2_n_89, sub_713_2_n_90, sub_713_2_n_91,
     sub_713_2_n_92, sub_713_2_n_93, sub_713_2_n_94, sub_713_2_n_95,
     sub_713_2_n_96, sub_713_2_n_97, sub_713_2_n_98, sub_713_2_n_99,
     sub_713_2_n_100, sub_713_2_n_101, sub_713_2_n_102, sub_713_2_n_103,
     sub_713_2_n_104, sub_713_2_n_105, sub_713_2_n_106, sub_713_2_n_107,
     sub_713_2_n_108, sub_713_2_n_109, sub_713_2_n_110, sub_713_2_n_111,
     sub_713_2_n_112, sub_713_2_n_113, sub_713_2_n_114, sub_713_2_n_115,
     sub_713_2_n_116, sub_713_2_n_117, sub_713_2_n_118, sub_713_2_n_119,
     sub_713_2_n_120, sub_713_2_n_121, sub_713_2_n_122, sub_713_2_n_123,
     sub_713_2_n_124, sub_713_2_n_125, sub_713_2_n_127, sub_713_2_n_128,
     sub_713_2_n_129, sub_713_2_n_130, sub_713_2_n_131, sub_713_2_n_132,
     sub_713_2_n_133, sub_713_2_n_135, sub_713_2_n_136, sub_713_2_n_138,
     sub_713_2_n_140, sub_713_2_n_141, sub_713_2_n_142, sub_713_2_n_145,
     sub_713_2_n_146, sub_713_2_n_149, sub_713_2_n_150, sub_713_2_n_151,
     sub_713_2_n_152, sub_713_2_n_156, sub_713_2_n_157, sub_713_2_n_158,
     sub_713_2_n_160, sub_713_2_n_161, sub_713_2_n_162, sub_713_2_n_163,
     sub_713_2_n_167, sub_713_2_n_168, sub_713_2_n_169, sub_713_2_n_174,
     sub_713_2_n_175, sub_713_2_n_176, sub_713_2_n_178, sub_713_2_n_186,
     sub_713_2_n_187, sub_713_2_n_188, sub_732_2_n_0, sub_732_2_n_1,
     sub_732_2_n_2, sub_732_2_n_3, sub_732_2_n_4, sub_732_2_n_5, sub_732_2_n_6,
     sub_732_2_n_7, sub_732_2_n_8, sub_732_2_n_9, sub_732_2_n_10, sub_732_2_n_11,
     sub_732_2_n_12, sub_732_2_n_13, sub_732_2_n_14, sub_732_2_n_15,
     sub_732_2_n_16, sub_732_2_n_17, sub_732_2_n_18, sub_732_2_n_19,
     sub_732_2_n_20, sub_732_2_n_21, sub_732_2_n_22, sub_732_2_n_23,
     sub_732_2_n_24, sub_732_2_n_25, sub_732_2_n_26, sub_732_2_n_27,
     sub_732_2_n_28, sub_732_2_n_29, sub_732_2_n_30, sub_732_2_n_31,
     sub_732_2_n_32, sub_732_2_n_33, sub_732_2_n_34, sub_732_2_n_35,
     sub_732_2_n_36, sub_732_2_n_37, sub_732_2_n_38, sub_732_2_n_39,
     sub_732_2_n_40, sub_732_2_n_41, sub_732_2_n_42, sub_732_2_n_43,
     sub_732_2_n_44, sub_732_2_n_45, sub_732_2_n_46, sub_732_2_n_47,
     sub_732_2_n_48, sub_732_2_n_49, sub_732_2_n_50, sub_732_2_n_51,
     sub_732_2_n_52, sub_732_2_n_53, sub_732_2_n_54, sub_732_2_n_55,
     sub_732_2_n_56, sub_732_2_n_57, sub_732_2_n_58, sub_732_2_n_59,
     sub_732_2_n_60, sub_732_2_n_61, sub_732_2_n_62, sub_732_2_n_63,
     sub_732_2_n_64, sub_732_2_n_65, sub_732_2_n_66, sub_732_2_n_67,
     sub_732_2_n_68, sub_732_2_n_69, sub_732_2_n_70, sub_732_2_n_71,
     sub_732_2_n_72, sub_732_2_n_73, sub_732_2_n_74, sub_732_2_n_75,
     sub_732_2_n_76, sub_732_2_n_78, sub_732_2_n_79, sub_732_2_n_80,
     sub_732_2_n_81, sub_732_2_n_82, sub_732_2_n_83, sub_732_2_n_84,
     sub_732_2_n_85, sub_732_2_n_86, sub_732_2_n_87, sub_732_2_n_88,
     sub_732_2_n_89, sub_732_2_n_90, sub_732_2_n_91, sub_732_2_n_92,
     sub_732_2_n_93, sub_732_2_n_94, sub_732_2_n_95, sub_732_2_n_96,
     sub_732_2_n_97, sub_732_2_n_98, sub_732_2_n_99, sub_732_2_n_100,
     sub_732_2_n_101, sub_732_2_n_102, sub_732_2_n_103, sub_732_2_n_104,
     sub_732_2_n_105, sub_732_2_n_106, sub_732_2_n_107, sub_732_2_n_108,
     sub_732_2_n_109, sub_732_2_n_110, sub_732_2_n_111, sub_732_2_n_112,
     sub_732_2_n_113, sub_732_2_n_114, sub_732_2_n_115, sub_732_2_n_116,
     sub_732_2_n_117, sub_732_2_n_118, sub_732_2_n_119, sub_732_2_n_120,
     sub_732_2_n_121, sub_732_2_n_122, sub_732_2_n_123, sub_732_2_n_124,
     sub_732_2_n_125, sub_732_2_n_126, sub_732_2_n_128, sub_732_2_n_129,
     sub_732_2_n_130, sub_732_2_n_131, sub_732_2_n_132, sub_732_2_n_133,
     sub_732_2_n_134, sub_732_2_n_135, sub_732_2_n_136, sub_732_2_n_138,
     sub_732_2_n_139, sub_732_2_n_140, sub_732_2_n_142, sub_732_2_n_144,
     sub_732_2_n_145, sub_732_2_n_146, sub_732_2_n_149, sub_732_2_n_150,
     sub_732_2_n_153, sub_732_2_n_154, sub_732_2_n_155, sub_732_2_n_156,
     sub_732_2_n_160, sub_732_2_n_161, sub_732_2_n_162, sub_732_2_n_164,
     sub_732_2_n_165, sub_732_2_n_166, sub_732_2_n_167, sub_732_2_n_168,
     sub_732_2_n_172, sub_732_2_n_173, sub_732_2_n_174, sub_732_2_n_179,
     sub_732_2_n_180, sub_732_2_n_181, sub_732_2_n_183, sub_732_2_n_191,
     sub_732_2_n_192, sub_732_2_n_193, sub_732_2_n_194, sub_751_2_n_0,
     sub_751_2_n_1, sub_751_2_n_2, sub_751_2_n_3, sub_751_2_n_4, sub_751_2_n_5,
     sub_751_2_n_6, sub_751_2_n_7, sub_751_2_n_8, sub_751_2_n_9, sub_751_2_n_10,
     sub_751_2_n_11, sub_751_2_n_12, sub_751_2_n_13, sub_751_2_n_14,
     sub_751_2_n_15, sub_751_2_n_16, sub_751_2_n_17, sub_751_2_n_18,
     sub_751_2_n_19, sub_751_2_n_20, sub_751_2_n_21, sub_751_2_n_22,
     sub_751_2_n_23, sub_751_2_n_24, sub_751_2_n_25, sub_751_2_n_26,
     sub_751_2_n_27, sub_751_2_n_28, sub_751_2_n_29, sub_751_2_n_30,
     sub_751_2_n_31, sub_751_2_n_32, sub_751_2_n_33, sub_751_2_n_34,
     sub_751_2_n_35, sub_751_2_n_36, sub_751_2_n_37, sub_751_2_n_38,
     sub_751_2_n_39, sub_751_2_n_40, sub_751_2_n_41, sub_751_2_n_42,
     sub_751_2_n_43, sub_751_2_n_44, sub_751_2_n_45, sub_751_2_n_46,
     sub_751_2_n_47, sub_751_2_n_48, sub_751_2_n_49, sub_751_2_n_50,
     sub_751_2_n_51, sub_751_2_n_52, sub_751_2_n_53, sub_751_2_n_54,
     sub_751_2_n_55, sub_751_2_n_56, sub_751_2_n_57, sub_751_2_n_58,
     sub_751_2_n_59, sub_751_2_n_60, sub_751_2_n_61, sub_751_2_n_62,
     sub_751_2_n_63, sub_751_2_n_64, sub_751_2_n_65, sub_751_2_n_66,
     sub_751_2_n_67, sub_751_2_n_68, sub_751_2_n_69, sub_751_2_n_70,
     sub_751_2_n_71, sub_751_2_n_72, sub_751_2_n_73, sub_751_2_n_74,
     sub_751_2_n_75, sub_751_2_n_76, sub_751_2_n_77, sub_751_2_n_79,
     sub_751_2_n_80, sub_751_2_n_81, sub_751_2_n_82, sub_751_2_n_83,
     sub_751_2_n_84, sub_751_2_n_85, sub_751_2_n_86, sub_751_2_n_87,
     sub_751_2_n_88, sub_751_2_n_89, sub_751_2_n_90, sub_751_2_n_91,
     sub_751_2_n_92, sub_751_2_n_93, sub_751_2_n_94, sub_751_2_n_95,
     sub_751_2_n_96, sub_751_2_n_97, sub_751_2_n_98, sub_751_2_n_99,
     sub_751_2_n_100, sub_751_2_n_101, sub_751_2_n_102, sub_751_2_n_103,
     sub_751_2_n_104, sub_751_2_n_105, sub_751_2_n_106, sub_751_2_n_107,
     sub_751_2_n_108, sub_751_2_n_109, sub_751_2_n_110, sub_751_2_n_111,
     sub_751_2_n_112, sub_751_2_n_113, sub_751_2_n_114, sub_751_2_n_115,
     sub_751_2_n_116, sub_751_2_n_117, sub_751_2_n_118, sub_751_2_n_119,
     sub_751_2_n_120, sub_751_2_n_121, sub_751_2_n_122, sub_751_2_n_123,
     sub_751_2_n_124, sub_751_2_n_125, sub_751_2_n_126, sub_751_2_n_127,
     sub_751_2_n_128, sub_751_2_n_129, sub_751_2_n_130, sub_751_2_n_131,
     sub_751_2_n_132, sub_751_2_n_134, sub_751_2_n_135, sub_751_2_n_137,
     sub_751_2_n_138, sub_751_2_n_139, sub_751_2_n_140, sub_751_2_n_142,
     sub_751_2_n_144, sub_751_2_n_145, sub_751_2_n_146, sub_751_2_n_149,
     sub_751_2_n_150, sub_751_2_n_153, sub_751_2_n_154, sub_751_2_n_155,
     sub_751_2_n_156, sub_751_2_n_160, sub_751_2_n_161, sub_751_2_n_162,
     sub_751_2_n_166, sub_751_2_n_167, sub_751_2_n_168, sub_751_2_n_172,
     sub_751_2_n_173, sub_751_2_n_178, sub_751_2_n_179, sub_751_2_n_180,
     sub_751_2_n_182, sub_751_2_n_183, sub_751_2_n_191, sub_751_2_n_192,
     sub_751_2_n_193, sub_751_2_n_194, sub_751_2_n_199, n_0, n_1, n_2, n_3, n_4,
     n_5, n_6, n_7, n_8, n_9, n_10, n_11, n_12, n_13, n_14, n_15, n_16, n_17,
     n_18, n_19, n_20, n_21, n_22, n_23, n_24, n_25, n_26, n_27, n_28, n_29,
     n_30, n_31, n_32, n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40, n_41,
     n_42, n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50, n_51, n_52, n_53,
     n_54, n_55, n_56, n_57, n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65,
     n_66, n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74, n_75, n_76, n_77,
     n_78, n_79, n_80, n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88, n_89,
     n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100, n_101,
     n_102, n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112,
     n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122, n_123,
     n_124, n_125, n_126, n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134,
     n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145,
     n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156,
     n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167,
     n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178,
     n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188, n_189,
     n_190, n_191, n_192, n_193, n_194, n_195, n_196, n_197, n_198, n_199, n_200,
     n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210, n_211,
     n_212, n_213, n_214, n_215, n_216, n_217, n_218, n_219, n_220, n_221, n_222,
     n_223, n_224, n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233,
     n_234, n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242, n_243, n_244,
     n_245, n_246, n_247, n_248, n_249, n_250, n_251, n_252, n_253, n_254, n_255,
     n_256, n_257, n_258, n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266,
     n_267, n_268, n_269, n_270, n_271, n_272, n_273, n_274, n_275, n_276, n_277,
     n_278, n_279, n_280, n_281, n_282, n_283, n_284, n_285, n_286, n_287, n_288,
     n_289, n_290, n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298, n_299,
     n_300, n_301, n_335, n_336, n_337, n_338, n_339, n_340, n_341, n_342, n_343,
     n_344, n_345, n_346, n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354,
     n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362, n_363, n_364, n_365,
     n_366, n_367, n_368, n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376,
     n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386, n_387,
     n_388, n_389, n_390, n_391, n_392, n_393, n_394, n_395, n_396, n_397, n_398,
     n_399, n_400, n_401, n_402, n_403, n_404, n_405, n_406, n_407, n_408, n_409,
     n_410, n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418, n_419, n_420,
     n_421, n_422, n_423, n_424, n_425, n_426, n_427, n_428, n_429, n_430, n_431,
     n_432, n_433, n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442,
     n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450, n_451, n_452, n_453,
     n_454, n_455, n_456, n_457, n_458, n_459, n_460, n_461, n_462, n_463, n_464,
     n_465, n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474, n_475,
     n_476, n_477, n_478, n_479, n_480, n_481, n_482, n_483, n_484, n_485, n_486,
     n_487, n_488, n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496, n_497,
     n_498, n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506, n_507, n_508,
     n_509, n_510, n_511, n_512, n_513, n_514, n_515, n_516, n_517, n_518, n_519,
     n_520, n_521, n_522, n_523, n_524, n_525, n_526, n_527, n_528, n_529, n_530,
     n_531, n_532, n_533, n_534, n_535, n_536, n_537, n_538, n_539, n_540, n_541,
     n_542, n_543, n_544, n_545, n_546, n_547, n_548, n_549, n_550, n_551, n_552,
     n_553, n_554, n_555, n_556, n_557, n_558, n_559, n_560, n_561, n_562, n_563,
     n_564, n_565, n_566, n_567, n_568, n_569, n_570, n_571, n_572, n_573, n_574,
     n_575, n_576, n_577, n_578, n_579, n_580, n_581, n_582, n_583, n_584, n_585,
     n_586, n_587, n_588, n_589, n_590, n_591, n_592, n_593, n_594, n_595, n_596,
     n_597, n_598, n_599, n_600, n_601, n_602, n_603, n_604, n_605, n_606, n_607,
     n_608, n_609, n_610, n_611, n_612, n_613, n_614, n_615, n_616, n_617, n_618,
     n_619, n_620, n_621, n_622, n_623, n_624, n_625, n_626, n_627, n_628, n_629,
     n_630, n_631, n_632, n_633, n_634, n_635, n_636, n_637, n_638, n_639, n_640,
     n_641, n_642, n_643, n_644, n_645, n_646, n_647, n_648, n_649, n_650, n_651,
     n_652, n_653, n_654, n_655, n_656, n_657, n_658, n_659, n_660, n_661, n_662,
     n_663, n_664, n_665, n_666, n_667, n_668, n_669, n_670, n_671, n_672, n_673,
     n_674, n_675, n_676, n_677, n_678, n_679, n_680, n_681, n_682, n_683, n_684,
     n_685, n_686, n_687, n_688, n_689, n_690, n_691, n_692, n_693, n_694, n_695,
     n_696, n_697, n_698, n_699, n_700, n_701, n_702, n_703, n_704, n_705, n_706,
     n_707, n_708, n_709, n_710, n_711, n_712, n_713, n_714, n_715, n_716, n_717,
     n_718, n_719, n_720, n_721, n_722, n_723, n_724, n_725, n_726, n_727, n_728,
     n_729, n_730, n_731, n_732, n_733, n_734, n_735, n_736, n_737, n_738, n_739,
     n_740, n_741, n_742, n_743, n_744, n_745, n_746, n_747, n_748, n_749, n_750,
     n_751, n_752, n_753, n_754, n_755, n_756, n_757, n_758, n_759, n_760, n_761,
     n_762, n_763, n_764, n_765, n_766, n_767, n_768, n_769, n_770, n_771, n_772,
     n_773, n_774, n_775, n_776, n_777, n_778, n_779, n_780, n_781, n_782, n_783,
     n_784, n_785, n_786, n_787, n_788, n_789, n_790, n_791, n_792, n_793, n_794,
     n_795, n_796, n_797, n_798, n_799, n_800, n_801, n_802, n_803, n_804, n_805,
     n_806, n_807, n_808, n_809, n_810, n_811, n_812, n_813, n_814, n_815, n_816,
     n_817, n_818, n_819, n_820, n_821, n_822, n_823, n_824, n_825, n_826, n_827,
     n_828, n_829, n_830, n_831, n_832, n_833, n_834, n_835, n_836, n_837, n_838,
     n_839, n_840, n_841, n_842, n_843, n_844, n_845, n_846, n_847, n_848, n_849,
     n_850, n_851, n_852, n_853, n_854, n_855, n_856, n_857, n_858, n_859, n_860,
     n_861, n_862, n_863, n_864, n_865, n_866, n_867, n_868, n_869, n_870, n_871,
     n_872, n_873, n_874, n_875, n_876, n_877, n_878, n_879, n_880, n_881, n_882,
     n_883, n_884, n_885, n_886, n_887, n_888, n_889, n_890, n_891, n_892, n_893,
     n_894, n_895, n_896, n_897, n_898, n_899, n_900, n_901, n_902, n_903, n_904,
     n_905, n_906, n_907, n_908, n_909, n_910, n_911, n_912, n_913, n_914, n_915,
     n_916, n_917, n_918, n_919, n_920, n_921, n_922, n_923, n_924, n_925, n_926,
     n_927, n_928, n_929, n_930, n_931, n_932, n_933, n_934, n_935, n_936, n_937,
     n_938, n_939, n_940, n_941, n_942, n_943, n_944, n_945, n_946, n_947, n_948,
     n_949, n_950, n_951, n_952, n_953, n_954, n_955, n_956, n_957, n_958, n_959,
     n_960, n_961, n_962, n_963, n_964, n_965, n_966, n_967, n_968, n_969, n_970,
     n_971, n_972, n_973, n_974, n_975, n_976, n_977, n_978, n_979, n_980, n_981,
     n_982, n_983, n_984, n_985, n_986, n_987, n_988, n_989, n_990, n_991, n_992,
     n_993, n_994, n_995, n_996, n_997, n_998, n_999, n_1000, n_1001, n_1002,
     n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011,
     n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020,
     n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029,
     n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038,
     n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047,
     n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056,
     n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065,
     n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074,
     n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083,
     n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092,
     n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101,
     n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110,
     n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119,
     n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128,
     n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137,
     n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146,
     n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155,
     n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164,
     n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173,
     n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182,
     n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191,
     n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200,
     n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209,
     n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218,
     n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227,
     n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236,
     n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245,
     n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254,
     n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263,
     n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272,
     n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281,
     n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290,
     n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299,
     n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308,
     n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317,
     n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326,
     n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335,
     n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344,
     n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353,
     n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362,
     n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371,
     n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380,
     n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389,
     n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398,
     n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, clk, clr, n_1441,
     n_1444, n_1445, n_1449, n_1450, n_1451, n_1456, n_1457, n_1458, n_1460,
     n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1473, n_1476, n_1477,
     n_1478, n_1479, n_1480, n_1481, n_1482, n_1489, n_1490, n_1491, n_1492,
     n_1493, n_1494, n_1496, n_1500, n_1502, n_1504, n_1505, n_1506, n_1507,
     n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1521, n_1522, n_1523,
     n_1524, n_1525, n_1526, n_1527, n_1528, n_1530, n_1531, n_1532, n_1533,
     n_1534, n_1535, n_1536, n_1537, n_1538, n_1540, n_1541, n_1542, n_1543,
     n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1561, n_1562,
     n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571,
     n_1572, n_1576, n_1579, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588,
     n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1599,
     n_1601, n_1607, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615,
     n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1636, n_1637,
     n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646,
     n_1647, n_1648, n_1649, n_1650, n_1652, n_1665, n_1666, n_1667, n_1668,
     n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677,
     n_1678, n_1679, n_1680, n_1688, n_1690, n_1692, n_1695, n_1696, n_1697,
     n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, n_1706,
     n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1725, n_1727, n_1728,
     n_1729, n_1730, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, n_1738,
     n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1764,
     n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773,
     n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782,
     n_1783, n_1788, n_1791, n_1799, n_1801, n_1802, n_1803, n_1804, n_1805,
     n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814,
     n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, n_1828, n_1841, n_1842,
     n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, n_1851,
     n_1852, n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860,
     n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, n_1889,
     n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896, n_1897, n_1898,
     n_1899, n_1900, n_1901, n_1902, n_1916, n_1921, n_1924, n_1925, n_1926,
     n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1934, n_1935, n_1936,
     n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1945,
     n_1946, n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, n_1976,
     n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, n_1985,
     n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992, n_2016, n_2017,
     n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, n_2025, n_2026,
     n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035,
     n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, n_2065, n_2067, n_2068,
     n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, n_2075, n_2076, n_2077,
     n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, n_2084, n_2085, n_2086,
     n_2087, n_2088, n_2089, n_2090, n_2105, n_2108, n_2116, n_2117, n_2118,
     n_2119, n_2120, n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, n_2127,
     n_2128, n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, n_2136,
     n_2137, n_2138, n_2139, n_2140, n_2141, n_2142, n_2160, n_2166, n_2169,
     n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, n_2178,
     n_2179, n_2180, n_2181, n_2182, n_2183, n_2184, n_2185, n_2186, n_2187,
     n_2188, n_2189, n_2190, n_2191, n_2192, n_2193, n_2194, n_2195, n_2196,
     n_2224, n_2225, n_2226, n_2227, n_2228, n_2229, n_2230, n_2231, n_2232,
     n_2233, n_2234, n_2235, n_2236, n_2237, n_2238, n_2239, n_2240, n_2241,
     n_2242, n_2243, n_2244, n_2245, n_2246, n_2247, n_2248, n_2249, n_2250,
     n_2251, n_2252, n_2254, n_2255, n_2256, n_2258, n_2259, n_2260, n_2282,
     n_2283, n_2284, n_2285, n_2286, n_2287, n_2288, n_2289, n_2290, n_2291,
     n_2292, n_2293, n_2294, n_2295, n_2296, n_2297, n_2298, n_2299, n_2300,
     n_2301, n_2302, n_2303, n_2304, n_2305, n_2306, n_2307, n_2308, n_2309,
     n_2310, n_2311, n_2312, n_2313, n_2314, n_2315, n_2316, n_2317, n_2318,
     n_2319, n_2320, n_2321, n_2322, n_2323, n_2324, n_2325, n_2326, n_2327,
     n_2328, n_2329, n_2330, n_2331, n_2332, n_2333, n_2334, n_2335, n_2336,
     n_2337, n_2338, n_2339, n_2340, n_2341, n_2342, n_2343, n_2344, n_2345,
     n_2346, n_2347, n_2348, n_2349, n_2350, n_2351, n_2352, n_2353, n_2354,
     n_2355, n_2356, n_2357, n_2358, n_2359, n_2360, n_2361, n_2362, n_2363,
     n_2364, n_2365, n_2366, n_2367, n_2368, n_2369, n_2370, n_2371, n_2372,
     n_2373, n_2374, n_2375, n_2376, n_2377, n_2378, n_2379, n_2380, n_2381,
     n_2382, n_2383, n_2384, n_2385, n_2386, n_2387, n_2388, n_2389, n_2390,
     n_2391, n_2392, n_2393, n_2394, n_2395, n_2396, n_2397, n_2398, n_2399,
     n_2400, n_2401, n_2402, n_2403, n_2404, n_2405, n_2406, n_2407, n_2408,
     n_2409, n_2410, n_2411, n_2412, n_2413, n_2414, n_2415, n_2416, n_2417,
     n_2418, n_2419, n_2420, n_2421, n_2422, n_2423, n_2424, n_2425, n_2426,
     n_2427, n_2428, n_2429, n_2430, n_2431, n_2432, n_2433, n_2434, n_2435,
     n_2436, n_2437, n_2438, n_2439, n_2440, n_2441, n_2442, n_2443, n_2444,
     n_2445, n_2446, n_2447, n_2448, n_2449, n_2450, n_2451, n_2452, n_2453,
     n_2454, n_2455, n_2456, n_2457, n_2458, n_2459, n_2460, n_2461, n_2462,
     n_2463, n_2464, n_2465, n_2466, n_2467, n_2468, n_2469, n_2470, n_2471,
     n_2472, n_2473, n_2474, n_2475, n_2476, n_2477, n_2478, n_2479, n_2480,
     n_2481, n_2482, n_2483, n_2484, n_2485, n_2486, n_2487, n_2488, n_2489,
     n_2490, n_2491, n_2492, n_2493, n_2494, n_2495, n_2496, n_2502, n_2503,
     n_2511, n_2516, n_2519, n_2520, n_2521, n_2522, n_2531, n_2532, n_2536,
     n_2542, n_2550, n_2551, n_2553, n_2554, n_2565, n_2567, n_2573, n_2576,
     n_2577, n_2578, n_2579, n_2580, n_2581, n_2582, n_2583, n_2590, n_2600,
     n_2602, n_2603, n_2607, n_2609, n_2618, n_2621, n_2622, n_2623, n_2624,
     n_2637, n_2652, n_2657, n_2658, n_2673, n_2674, n_2677, n_2678, n_2682,
     n_2694, n_2695, n_2696, n_2698, n_2717, n_2719, n_2736, n_2737, n_2738,
     n_2744, n_2747, n_2748, n_2749, n_2753, n_2775, n_2781, n_2805, n_2826,
     n_2829, n_2833, n_2863, n_2889, n_2897, n_2944, n_2947, n_2949, n_2972,
     n_2978, n_2979, n_3009, n_3030, n_3034, n_3036, n_3038, n_3042, n_3043,
     n_3044, n_3045, n_3047, n_3048, n_3049, n_3050, n_3051, n_3052, n_3053,
     n_3054, n_3055, n_3056, n_3057, n_3058, n_3059, n_3060, n_3061, n_3062,
     n_3063, n_3064, n_3065, n_3066, n_3067, n_3068, n_3069, n_3070, n_3071,
     n_3072, n_3080, n_3083, n_3092, n_3095, n_3099, n_3102, n_3105, n_3106,
     n_3109, n_3113, n_3117, n_3118, n_3119, n_3121, n_3122, n_3123, n_3124,
     n_3125, n_3126, n_3127, n_3128, n_3129, n_3131, n_3134, n_3136, n_3137,
     n_3138, n_3139, n_3140, n_3141, n_3142, n_3143, n_3144, n_3145, n_3146,
     n_3147, n_3148, n_3149, n_3150, n_3152, n_3153, n_3154, n_3159, n_3161,
     n_3164, n_3165, n_3166, n_3167, n_3169, n_3170, n_3171, n_3172, n_3173,
     n_3174, n_3175, n_3176, n_3177, n_3178, n_3179, n_3180, n_3181, n_3182,
     n_3183, n_3185, n_3188, n_3189, n_3190, n_2606, n_3192, n_3193, n_3194,
     n_3197, n_3199, n_3200, n_3201, n_3202, n_3204, n_3205, n_3207, n_3208,
     n_3209, n_3210, n_3211, n_3212, n_3213, n_3214, n_3215, n_3216, n_3217,
     n_3218, n_3219, n_3220, n_3221, n_3222, n_3223, n_3224, n_3225, n_3226,
     n_3227, n_3228, n_3229, n_3230, n_3231, n_3232, n_3233, n_3234, n_3235,
     n_3236, n_3237, n_3238, n_3239, n_3240, n_3241, n_3242, n_3243, n_3244,
     n_3245, n_3246, n_3247, n_3248, n_3249, n_3250, n_3251, n_3252, n_3253,
     n_3254, n_3255, n_3256, n_3257, n_3258, n_3259, n_3260, n_3261, n_3262,
     n_3263, n_3264, n_3265, n_3266, n_3267, n_3268, n_3269, n_3270, n_3271,
     n_3272, n_3273, n_3274, n_3275, n_3276, n_3277, n_3278, n_3279, n_3280,
     n_3281, n_3282, n_3283, n_3284, n_3285, n_3286, n_3287, n_3288, n_3289,
     n_3290, n_3291, n_3292, n_3293, n_3294, n_3295, n_3296, n_3297, n_3298,
     n_3299, n_3300, n_3301, n_3302, n_3303, n_3304, n_3305, n_3306, n_3307,
     n_3308, n_3309, n_3312, n_3314, n_3316, n_3317, n_3318, n_3319, n_3320,
     n_3321, n_3322, n_3323, n_3324, n_3325, n_3326, n_3327, n_3328, n_3329,
     n_3330, n_3331, n_3332, n_3333, n_3337, n_3338, n_3339, n_3341, n_3343,
     n_3344, n_3345, n_3346, n_3347, n_3348, n_3349, n_3350, n_3351, n_3352,
     n_3353, n_3354, n_3355, n_3356, n_3357, n_3358, n_3359, n_3360, n_3361,
     n_3362, n_3363, n_3364, n_3365, n_3366, n_3367, n_3368, n_3369, n_3370,
     n_3371, n_3372, n_3373, n_3374, n_3375, n_3376, n_3377, n_3378, n_3379,
     n_3380, n_3381, n_3382, n_3383, n_3384, n_3385, n_3386, n_3387, n_3388,
     n_3389, n_3390, n_3391, n_3392, n_3393, n_3394, n_3395, n_3396, n_3397,
     n_3398, n_3399, n_3400, n_3401, n_3402, n_3403, n_3404, n_3405, n_3406,
     n_3407, n_3408, n_3409, n_3410, n_3411, n_3412, n_3413, n_3414, n_3415,
     n_3416, n_3417, n_3418, n_3419, n_3420, n_3421, n_3422, n_3423, n_3424,
     n_3425, n_3426, n_3427, n_3428, n_3429, n_3430, n_3431, n_3432, n_3433,
     n_3434, n_3435, n_3436, n_3437, n_3438, n_3439, n_3440, n_3441, n_3442,
     n_3443, n_3444, n_3445, n_3446, n_3447, n_3448, n_3449, n_3450, n_3451,
     n_3452, n_3453, n_3454, n_3455, n_3456, n_3457, n_3458, n_3459, n_3460,
     n_3461, n_3462, n_3463, n_3464, n_3465, n_3466, n_3467, n_3468, n_3469,
     n_3470, n_3471, n_3472, n_3473, n_3474, n_3475, n_3476, n_3477, n_3478,
     n_3479, n_3480, n_3481, n_3482, n_3483, n_3484, n_3485, n_3486, n_3487,
     n_3488, n_3489, n_3490, n_3491, n_3492, n_3493, n_3494, n_3495, n_3496,
     n_3497, n_3498, n_3499, n_3500, n_3501, n_3502, n_3503, n_3504, n_3505,
     n_3506, n_3507, n_3508, n_3509, n_3510, n_3511, n_3512, n_3513, n_3514,
     n_3515, n_3516, n_3517, n_3518, n_3519, n_3520, n_3521, n_3522, n_3523,
     n_3524, n_3525, n_3526, n_3527, n_3528, n_3529, n_3530, n_3531, n_3532,
     n_3533, n_3534, n_3535, n_3536, n_3537, n_3538, n_3540, n_3541, n_3542,
     n_3543, n_3544, n_3545, n_3546, n_3547, n_3548, n_3549, n_3550, n_3551,
     n_3552, n_3553, n_3554, n_3555, n_3556, n_3557, n_3558, n_3559, n_3560,
     n_3561, n_3562, n_3563, n_3564, n_3565, n_3566, n_3567, n_3568, n_3569,
     n_3570, n_3571, n_3572, n_3573, n_3574, n_3575, n_3576, n_3577, n_3578,
     n_3579, n_3580, n_3581, n_3582, n_3583, n_3584, n_3585, n_3586, n_3587,
     n_3588, n_3589, n_3591, n_3592, n_3593, n_3594, n_3595, n_3596, n_3597,
     n_3598, n_3599, n_3600, n_3601, n_3602, n_3603, n_3604, n_3605, n_3606,
     n_3607, n_3608, n_3609, n_3610, n_3611, n_3612, n_3613, n_3614, n_3615,
     n_3616, n_3617, n_3618, n_3619, n_3620, n_3621, n_3622, n_3623, n_3624,
     n_3625, n_3626, n_3627, n_3628, n_3629, n_3630, n_3631, n_3632, n_3633,
     n_3634, n_3635, n_3636, n_3637, n_3638, n_3639, n_3640, n_3641, n_3642,
     n_3643, n_3644, n_3645, n_3646, n_3647, n_3648, n_3649, n_3650, n_3651,
     n_3652, n_3653, n_3654, n_3655, n_3656, n_3657, n_3658, n_3659, n_3660,
     n_3661, n_3662, n_3663, n_3664, n_3665, n_3666, n_3667, n_3668, n_3669,
     n_3670, n_3671, n_3672, n_3673, n_3674, n_3675, n_3676, n_3677, n_3678,
     n_3679, n_3680, n_3681, n_3682, n_3683, n_3684, n_3685, n_3686, n_3687,
     n_3688, n_3689, n_3690, n_3692, n_3693, n_3694, n_3695, n_3696, n_3697,
     n_3699, n_3700, n_3701, n_3702, n_3703, n_3704, n_3705, n_3706, n_3707,
     n_3708, n_3709, n_3710, n_3711, n_3712, n_3713, n_3714, n_3715, n_3716,
     n_3717, n_3718, n_3719, n_3720, n_3721, n_3722, n_3723, n_3724, n_3725,
     n_3726, n_3727, n_3728, n_3729, n_3730, n_3731, n_3732, n_3733, n_3734,
     n_3735, n_3736, n_3737, n_3738, n_3739, n_3740, n_3741, n_3742, n_3743,
     n_3744, n_3745, n_3746, n_3747, n_3748, n_3749, in2_95_0_, in2_95_1_,
     in2_95_2_, in2_95_3_, in2_95_4_, in2_95_5_, in2_95_6_, in2_95_7_, in2_95_8_,
     in2_95_9_, in2_95_10_, in2_95_11_, in2_95_12_, in2_95_13_, in2_95_14_,
     in2_95_15_, in2_95_16_, in2_95_17_, in2_95_18_, in2_95_19_, in2_95_20_,
     in2_95_21_, in2_95_22_, in2_95_23_, in2_95_24_, in2_95_25_, in2_95_26_,
     in2_95_27_, in2_95_28_, in2_95_29_, in2_95_30_, in2_95_31_, in;
assign n_1405 = in2_95_31_;
assign n_1373 = n_1405;
assign n_1341 = n_1373;
assign n_1309 = n_1341;
assign n_1277 = n_1309;
assign n_1245 = n_1277;
assign n_1213 = n_1245;
assign n_1181 = n_1213;
assign n_1149 = n_1181;
assign {out1[31]} = n_1149;
assign n_1404 = in2_95_30_;
assign n_1372 = n_1404;
assign n_1340 = n_1372;
assign n_1308 = n_1340;
assign n_1276 = n_1308;
assign n_1244 = n_1276;
assign n_1212 = n_1244;
assign n_1180 = n_1212;
assign n_1148 = n_1180;
assign {out1[30]} = n_1148;
assign n_1403 = in2_95_29_;
assign n_1371 = n_1403;
assign n_1339 = n_1371;
assign n_1307 = n_1339;
assign n_1275 = n_1307;
assign n_1243 = n_1275;
assign n_1211 = n_1243;
assign n_1179 = n_1211;
assign n_1147 = n_1179;
assign {out1[29]} = n_1147;
assign n_1402 = in2_95_28_;
assign n_1370 = n_1402;
assign n_1338 = n_1370;
assign n_1306 = n_1338;
assign n_1274 = n_1306;
assign n_1242 = n_1274;
assign n_1210 = n_1242;
assign n_1178 = n_1210;
assign n_1146 = n_1178;
assign {out1[28]} = n_1146;
assign n_1401 = in2_95_27_;
assign n_1369 = n_1401;
assign n_1337 = n_1369;
assign n_1305 = n_1337;
assign n_1273 = n_1305;
assign n_1241 = n_1273;
assign n_1209 = n_1241;
assign n_1177 = n_1209;
assign n_1145 = n_1177;
assign {out1[27]} = n_1145;
assign n_1400 = in2_95_26_;
assign n_1368 = n_1400;
assign n_1336 = n_1368;
assign n_1304 = n_1336;
assign n_1272 = n_1304;
assign n_1240 = n_1272;
assign n_1208 = n_1240;
assign n_1176 = n_1208;
assign n_1144 = n_1176;
assign {out1[26]} = n_1144;
assign n_1399 = in2_95_25_;
assign n_1367 = n_1399;
assign n_1335 = n_1367;
assign n_1303 = n_1335;
assign n_1271 = n_1303;
assign n_1239 = n_1271;
assign n_1207 = n_1239;
assign n_1175 = n_1207;
assign n_1143 = n_1175;
assign {out1[25]} = n_1143;
assign n_1398 = in2_95_24_;
assign n_1366 = n_1398;
assign n_1334 = n_1366;
assign n_1302 = n_1334;
assign n_1270 = n_1302;
assign n_1238 = n_1270;
assign n_1206 = n_1238;
assign n_1174 = n_1206;
assign n_1142 = n_1174;
assign {out1[24]} = n_1142;
assign n_1397 = in2_95_23_;
assign n_1365 = n_1397;
assign n_1333 = n_1365;
assign n_1301 = n_1333;
assign n_1269 = n_1301;
assign n_1237 = n_1269;
assign n_1205 = n_1237;
assign n_1173 = n_1205;
assign n_1141 = n_1173;
assign {out1[23]} = n_1141;
assign n_1396 = in2_95_22_;
assign n_1364 = n_1396;
assign n_1332 = n_1364;
assign n_1300 = n_1332;
assign n_1268 = n_1300;
assign n_1236 = n_1268;
assign n_1204 = n_1236;
assign n_1172 = n_1204;
assign n_1140 = n_1172;
assign {out1[22]} = n_1140;
assign n_1395 = in2_95_21_;
assign n_1363 = n_1395;
assign n_1331 = n_1363;
assign n_1299 = n_1331;
assign n_1267 = n_1299;
assign n_1235 = n_1267;
assign n_1203 = n_1235;
assign n_1171 = n_1203;
assign n_1139 = n_1171;
assign {out1[21]} = n_1139;
assign n_1394 = in2_95_20_;
assign n_1362 = n_1394;
assign n_1330 = n_1362;
assign n_1298 = n_1330;
assign n_1266 = n_1298;
assign n_1234 = n_1266;
assign n_1202 = n_1234;
assign n_1170 = n_1202;
assign n_1138 = n_1170;
assign {out1[20]} = n_1138;
assign n_1393 = in2_95_19_;
assign n_1361 = n_1393;
assign n_1329 = n_1361;
assign n_1297 = n_1329;
assign n_1265 = n_1297;
assign n_1233 = n_1265;
assign n_1201 = n_1233;
assign n_1169 = n_1201;
assign n_1137 = n_1169;
assign {out1[19]} = n_1137;
assign n_1392 = in2_95_18_;
assign n_1360 = n_1392;
assign n_1328 = n_1360;
assign n_1296 = n_1328;
assign n_1264 = n_1296;
assign n_1232 = n_1264;
assign n_1200 = n_1232;
assign n_1168 = n_1200;
assign n_1136 = n_1168;
assign {out1[18]} = n_1136;
assign n_1391 = in2_95_17_;
assign n_1359 = n_1391;
assign n_1327 = n_1359;
assign n_1295 = n_1327;
assign n_1263 = n_1295;
assign n_1231 = n_1263;
assign n_1199 = n_1231;
assign n_1167 = n_1199;
assign n_1135 = n_1167;
assign {out1[17]} = n_1135;
assign n_1390 = in2_95_16_;
assign n_1358 = n_1390;
assign n_1326 = n_1358;
assign n_1294 = n_1326;
assign n_1262 = n_1294;
assign n_1230 = n_1262;
assign n_1198 = n_1230;
assign n_1166 = n_1198;
assign n_1134 = n_1166;
assign {out1[16]} = n_1134;
assign n_1389 = in2_95_15_;
assign n_1357 = n_1389;
assign n_1325 = n_1357;
assign n_1293 = n_1325;
assign n_1261 = n_1293;
assign n_1229 = n_1261;
assign n_1197 = n_1229;
assign n_1165 = n_1197;
assign n_1133 = n_1165;
assign {out1[15]} = n_1133;
assign n_1388 = in2_95_14_;
assign n_1356 = n_1388;
assign n_1324 = n_1356;
assign n_1292 = n_1324;
assign n_1260 = n_1292;
assign n_1228 = n_1260;
assign n_1196 = n_1228;
assign n_1164 = n_1196;
assign n_1132 = n_1164;
assign {out1[14]} = n_1132;
assign n_1387 = in2_95_13_;
assign n_1355 = n_1387;
assign n_1323 = n_1355;
assign n_1291 = n_1323;
assign n_1259 = n_1291;
assign n_1227 = n_1259;
assign n_1195 = n_1227;
assign n_1163 = n_1195;
assign n_1131 = n_1163;
assign {out1[13]} = n_1131;
assign n_1386 = in2_95_12_;
assign n_1354 = n_1386;
assign n_1322 = n_1354;
assign n_1290 = n_1322;
assign n_1258 = n_1290;
assign n_1226 = n_1258;
assign n_1194 = n_1226;
assign n_1162 = n_1194;
assign n_1130 = n_1162;
assign {out1[12]} = n_1130;
assign n_1385 = in2_95_11_;
assign n_1353 = n_1385;
assign n_1321 = n_1353;
assign n_1289 = n_1321;
assign n_1257 = n_1289;
assign n_1225 = n_1257;
assign n_1193 = n_1225;
assign n_1161 = n_1193;
assign n_1129 = n_1161;
assign {out1[11]} = n_1129;
assign n_1384 = in2_95_10_;
assign n_1352 = n_1384;
assign n_1320 = n_1352;
assign n_1288 = n_1320;
assign n_1256 = n_1288;
assign n_1224 = n_1256;
assign n_1192 = n_1224;
assign n_1160 = n_1192;
assign n_1128 = n_1160;
assign {out1[10]} = n_1128;
assign n_1383 = in2_95_9_;
assign n_1351 = n_1383;
assign n_1319 = n_1351;
assign n_1287 = n_1319;
assign n_1255 = n_1287;
assign n_1223 = n_1255;
assign n_1191 = n_1223;
assign n_1159 = n_1191;
assign n_1127 = n_1159;
assign {out1[9]} = n_1127;
assign n_1382 = in2_95_8_;
assign n_1350 = n_1382;
assign n_1318 = n_1350;
assign n_1286 = n_1318;
assign n_1254 = n_1286;
assign n_1222 = n_1254;
assign n_1190 = n_1222;
assign n_1158 = n_1190;
assign n_1126 = n_1158;
assign {out1[8]} = n_1126;
assign n_1381 = in2_95_7_;
assign n_1349 = n_1381;
assign n_1317 = n_1349;
assign n_1285 = n_1317;
assign n_1253 = n_1285;
assign n_1221 = n_1253;
assign n_1189 = n_1221;
assign n_1157 = n_1189;
assign n_1125 = n_1157;
assign {out1[7]} = n_1125;
assign n_1380 = in2_95_6_;
assign n_1348 = n_1380;
assign n_1316 = n_1348;
assign n_1284 = n_1316;
assign n_1252 = n_1284;
assign n_1220 = n_1252;
assign n_1188 = n_1220;
assign n_1156 = n_1188;
assign n_1124 = n_1156;
assign {out1[6]} = n_1124;
assign n_1379 = in2_95_5_;
assign n_1347 = n_1379;
assign n_1315 = n_1347;
assign n_1283 = n_1315;
assign n_1251 = n_1283;
assign n_1219 = n_1251;
assign n_1187 = n_1219;
assign n_1155 = n_1187;
assign n_1123 = n_1155;
assign {out1[5]} = n_1123;
assign n_1378 = in2_95_4_;
assign n_1346 = n_1378;
assign n_1314 = n_1346;
assign n_1282 = n_1314;
assign n_1250 = n_1282;
assign n_1218 = n_1250;
assign n_1186 = n_1218;
assign n_1154 = n_1186;
assign n_1122 = n_1154;
assign {out1[4]} = n_1122;
assign n_1377 = in2_95_3_;
assign n_1345 = n_1377;
assign n_1313 = n_1345;
assign n_1281 = n_1313;
assign n_1249 = n_1281;
assign n_1217 = n_1249;
assign n_1185 = n_1217;
assign n_1153 = n_1185;
assign n_1121 = n_1153;
assign {out1[3]} = n_1121;
assign n_1376 = in2_95_2_;
assign n_1344 = n_1376;
assign n_1312 = n_1344;
assign n_1280 = n_1312;
assign n_1248 = n_1280;
assign n_1216 = n_1248;
assign n_1184 = n_1216;
assign n_1152 = n_1184;
assign n_1120 = n_1152;
assign {out1[2]} = n_1120;
assign n_1375 = in2_95_1_;
assign n_1343 = n_1375;
assign n_1311 = n_1343;
assign n_1279 = n_1311;
assign n_1247 = n_1279;
assign n_1215 = n_1247;
assign n_1183 = n_1215;
assign n_1151 = n_1183;
assign n_1119 = n_1151;
assign {out1[1]} = n_1119;
assign n_1374 = in2_95_0_;
assign n_1342 = n_1374;
assign n_1310 = n_1342;
assign n_1278 = n_1310;
assign n_1246 = n_1278;
assign n_1214 = n_1246;
assign n_1182 = n_1214;
assign n_1150 = n_1182;
assign n_1118 = n_1150;
assign {out1[0]} = n_1118;
 reg retime_s1_3_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_3_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_3_reg_reg_IQ <= {in1[24]};
     end
 assign n_1115 = retime_s1_3_reg_reg_IQ;
 reg retime_s1_4_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_4_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_4_reg_reg_IQ <= {in2[25]};
     end
 assign n_726 = retime_s1_4_reg_reg_IQ;
 reg retime_s1_5_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_5_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_5_reg_reg_IQ <= n_1496;
     end
 assign n_725 = retime_s1_5_reg_reg_IQ;
 reg retime_s1_6_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_6_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_6_reg_reg_IQ <= n_3231;
     end
 assign n_724 = retime_s1_6_reg_reg_IQ;
 reg retime_s1_9_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_9_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_9_reg_reg_IQ <= n_1480;
     end
 assign n_721 = retime_s1_9_reg_reg_IQ;
 reg retime_s1_12_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_12_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_12_reg_reg_IQ <= n_1479;
     end
 assign n_718 = retime_s1_12_reg_reg_IQ;
 reg retime_s1_17_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_17_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_17_reg_reg_IQ <= {in2[23]};
     end
 assign n_713 = retime_s1_17_reg_reg_IQ;
 reg retime_s1_18_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_18_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_18_reg_reg_IQ <= n_1530;
     end
 assign n_712 = retime_s1_18_reg_reg_IQ;
 reg retime_s1_19_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_19_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_19_reg_reg_IQ <= n_3230;
     end
 assign n_711 = retime_s1_19_reg_reg_IQ;
 reg retime_s1_22_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_22_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_22_reg_reg_IQ <= sub_257_2_n_49;
     end
 assign n_708 = retime_s1_22_reg_reg_IQ;
 reg retime_s1_23_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_23_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_23_reg_reg_IQ <= sub_257_2_n_33;
     end
 assign n_707 = retime_s1_23_reg_reg_IQ;
 reg retime_s1_25_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_25_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_25_reg_reg_IQ <= {in1[4]};
     end
 assign n_705 = retime_s1_25_reg_reg_IQ;
 reg retime_s1_26_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_26_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_26_reg_reg_IQ <= sub_257_2_n_48;
     end
 assign n_695 = retime_s1_26_reg_reg_IQ;
 reg retime_s1_27_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_27_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_27_reg_reg_IQ <= n_1478;
     end
 assign n_694 = retime_s1_27_reg_reg_IQ;
 reg retime_s1_28_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_28_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_28_reg_reg_IQ <= {in1[12]};
     end
 assign n_693 = retime_s1_28_reg_reg_IQ;
 reg retime_s1_29_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_29_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_29_reg_reg_IQ <= {in1[7]};
     end
 assign n_683 = retime_s1_29_reg_reg_IQ;
 reg retime_s1_33_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_33_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_33_reg_reg_IQ <= {in1[26]};
     end
 assign n_670 = retime_s1_33_reg_reg_IQ;
 reg retime_s1_34_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_34_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_34_reg_reg_IQ <= {in1[6]};
     end
 assign n_660 = retime_s1_34_reg_reg_IQ;
 reg retime_s1_36_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_36_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_36_reg_reg_IQ <= n_3225;
     end
 assign n_649 = retime_s1_36_reg_reg_IQ;
 reg retime_s1_37_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_37_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_37_reg_reg_IQ <= n_3226;
     end
 assign n_648 = retime_s1_37_reg_reg_IQ;
 reg retime_s1_38_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_38_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_38_reg_reg_IQ <= n_1481;
     end
 assign n_647 = retime_s1_38_reg_reg_IQ;
 reg retime_s1_39_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_39_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_39_reg_reg_IQ <= n_1473;
     end
 assign n_646 = retime_s1_39_reg_reg_IQ;
 reg retime_s1_40_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_40_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_40_reg_reg_IQ <= sub_314_2_n_18;
     end
 assign n_645 = retime_s1_40_reg_reg_IQ;
 reg retime_s1_41_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_41_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_41_reg_reg_IQ <= sub_276_2_n_16;
     end
 assign n_644 = retime_s1_41_reg_reg_IQ;
 reg retime_s1_42_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_42_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_42_reg_reg_IQ <= {in2[26]};
     end
 assign n_643 = retime_s1_42_reg_reg_IQ;
 reg retime_s1_43_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_43_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_43_reg_reg_IQ <= {in1[5]};
     end
 assign n_642 = retime_s1_43_reg_reg_IQ;
 reg retime_s1_48_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_48_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_48_reg_reg_IQ <= {in1[28]};
     end
 assign n_628 = retime_s1_48_reg_reg_IQ;
 reg retime_s1_50_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_50_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_50_reg_reg_IQ <= n_1482;
     end
 assign n_617 = retime_s1_50_reg_reg_IQ;
 reg retime_s1_53_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_53_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_53_reg_reg_IQ <= {in1[18]};
     end
 assign n_614 = retime_s1_53_reg_reg_IQ;
 reg retime_s1_54_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_54_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_54_reg_reg_IQ <= {in1[21]};
     end
 assign n_604 = retime_s1_54_reg_reg_IQ;
 reg retime_s1_55_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_55_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_55_reg_reg_IQ <= {in1[29]};
     end
 assign n_594 = retime_s1_55_reg_reg_IQ;
 reg retime_s1_63_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_63_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_63_reg_reg_IQ <= n_1550;
     end
 assign n_285 = retime_s1_63_reg_reg_IQ;
 reg retime_s1_64_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_64_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_64_reg_reg_IQ <= sub_333_2_n_18;
     end
 assign n_576 = retime_s1_64_reg_reg_IQ;
 reg retime_s1_72_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_72_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_72_reg_reg_IQ <= {in1[17]};
     end
 assign n_568 = retime_s1_72_reg_reg_IQ;
 reg retime_s1_73_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_73_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_73_reg_reg_IQ <= {in1[27]};
     end
 assign n_558 = retime_s1_73_reg_reg_IQ;
 reg retime_s1_74_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_74_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_74_reg_reg_IQ <= {in1[25]};
     end
 assign n_548 = retime_s1_74_reg_reg_IQ;
 reg retime_s1_75_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_75_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_75_reg_reg_IQ <= {in1[3]};
     end
 assign n_538 = retime_s1_75_reg_reg_IQ;
 reg retime_s1_76_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_76_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_76_reg_reg_IQ <= sub_257_2_n_39;
     end
 assign n_528 = retime_s1_76_reg_reg_IQ;
 reg retime_s1_77_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_77_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_77_reg_reg_IQ <= {in1[15]};
     end
 assign n_527 = retime_s1_77_reg_reg_IQ;
 reg retime_s1_88_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_88_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_88_reg_reg_IQ <= {in1[31]};
     end
 assign n_507 = retime_s1_88_reg_reg_IQ;
 reg retime_s1_92_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_92_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_92_reg_reg_IQ <= n_3164;
     end
 assign n_494 = retime_s1_92_reg_reg_IQ;
 reg retime_s1_97_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_97_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_97_reg_reg_IQ <= {in2[24]};
     end
 assign n_489 = retime_s1_97_reg_reg_IQ;
 reg retime_s1_98_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_98_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_98_reg_reg_IQ <= n_1512;
     end
 assign n_488 = retime_s1_98_reg_reg_IQ;
 reg retime_s1_99_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_99_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_99_reg_reg_IQ <= sub_295_2_n_19;
     end
 assign n_487 = retime_s1_99_reg_reg_IQ;
 reg retime_s1_100_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_100_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_100_reg_reg_IQ <= {in1[20]};
     end
 assign n_486 = retime_s1_100_reg_reg_IQ;
 reg retime_s1_101_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_101_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_101_reg_reg_IQ <= {in1[16]};
     end
 assign n_476 = retime_s1_101_reg_reg_IQ;
 reg retime_s1_102_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_102_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_102_reg_reg_IQ <= {in1[23]};
     end
 assign n_466 = retime_s1_102_reg_reg_IQ;
 reg retime_s1_103_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_103_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_103_reg_reg_IQ <= {in1[19]};
     end
 assign n_456 = retime_s1_103_reg_reg_IQ;
 reg retime_s1_105_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_105_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_105_reg_reg_IQ <= {in1[8]};
     end
 assign n_445 = retime_s1_105_reg_reg_IQ;
 reg retime_s1_106_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_106_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_106_reg_reg_IQ <= {in1[11]};
     end
 assign n_435 = retime_s1_106_reg_reg_IQ;
 reg retime_s1_107_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_107_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_107_reg_reg_IQ <= {in1[2]};
     end
 assign n_425 = retime_s1_107_reg_reg_IQ;
 reg retime_s1_108_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_108_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_108_reg_reg_IQ <= {in1[30]};
     end
 assign n_415 = retime_s1_108_reg_reg_IQ;
 reg retime_s1_113_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_113_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_113_reg_reg_IQ <= {in1[9]};
     end
 assign n_401 = retime_s1_113_reg_reg_IQ;
 reg retime_s1_114_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_114_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_114_reg_reg_IQ <= {in1[1]};
     end
 assign n_391 = retime_s1_114_reg_reg_IQ;
 reg retime_s1_120_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_120_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_120_reg_reg_IQ <= {in1[14]};
     end
 assign n_376 = retime_s1_120_reg_reg_IQ;
 reg retime_s1_122_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_122_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_122_reg_reg_IQ <= {in1[10]};
     end
 assign n_365 = retime_s1_122_reg_reg_IQ;
 reg retime_s1_123_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_123_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_123_reg_reg_IQ <= {in1[13]};
     end
 assign n_355 = retime_s1_123_reg_reg_IQ;
 reg retime_s1_125_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_125_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_125_reg_reg_IQ <= {in1[22]};
     end
 assign n_344 = retime_s1_125_reg_reg_IQ;
 reg retime_s2_3_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_3_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_3_reg_reg_IQ <= n_1115;
     end
 assign n_1114 = retime_s2_3_reg_reg_IQ;
 reg retime_s2_4_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_4_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_4_reg_reg_IQ <= n_1534;
     end
 assign n_750 = retime_s2_4_reg_reg_IQ;
 reg retime_s2_5_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_5_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_5_reg_reg_IQ <= n_1537;
     end
 assign n_749 = retime_s2_5_reg_reg_IQ;
 reg retime_s2_6_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_6_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_6_reg_reg_IQ <= sub_333_2_n_3;
     end
 assign n_748 = retime_s2_6_reg_reg_IQ;
 reg retime_s2_7_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_7_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_7_reg_reg_IQ <= n_1538;
     end
 assign n_747 = retime_s2_7_reg_reg_IQ;
 reg retime_s2_8_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_8_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_8_reg_reg_IQ <= sub_333_2_n_35;
     end
 assign n_746 = retime_s2_8_reg_reg_IQ;
 reg retime_s2_9_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_9_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_9_reg_reg_IQ <= sub_333_2_n_62;
     end
 assign n_745 = retime_s2_9_reg_reg_IQ;
 reg retime_s2_10_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_10_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_10_reg_reg_IQ <= sub_333_2_n_20;
     end
 assign n_744 = retime_s2_10_reg_reg_IQ;
 reg retime_s2_11_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_11_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_11_reg_reg_IQ <= n_1532;
     end
 assign n_743 = retime_s2_11_reg_reg_IQ;
 reg retime_s2_12_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_12_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_12_reg_reg_IQ <= n_1535;
     end
 assign n_742 = retime_s2_12_reg_reg_IQ;
 reg retime_s2_13_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_13_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_13_reg_reg_IQ <= sub_333_2_n_46;
     end
 assign n_741 = retime_s2_13_reg_reg_IQ;
 reg retime_s2_14_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_14_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_14_reg_reg_IQ <= sub_333_2_n_39;
     end
 assign n_740 = retime_s2_14_reg_reg_IQ;
 reg retime_s2_15_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_15_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_15_reg_reg_IQ <= sub_333_2_n_44;
     end
 assign n_739 = retime_s2_15_reg_reg_IQ;
 reg retime_s2_16_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_16_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_16_reg_reg_IQ <= n_1533;
     end
 assign n_738 = retime_s2_16_reg_reg_IQ;
 reg retime_s2_17_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_17_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_17_reg_reg_IQ <= n_3044;
     end
 assign n_737 = retime_s2_17_reg_reg_IQ;
 reg retime_s2_18_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_18_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_18_reg_reg_IQ <= sub_333_2_n_29;
     end
 assign n_736 = retime_s2_18_reg_reg_IQ;
 reg retime_s2_19_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_19_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_19_reg_reg_IQ <= n_1549;
     end
 assign n_735 = retime_s2_19_reg_reg_IQ;
 reg retime_s2_20_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_20_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_20_reg_reg_IQ <= n_1536;
     end
 assign n_734 = retime_s2_20_reg_reg_IQ;
 reg retime_s2_21_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_21_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_21_reg_reg_IQ <= sub_333_2_n_1;
     end
 assign n_733 = retime_s2_21_reg_reg_IQ;
 reg retime_s2_22_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_22_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_22_reg_reg_IQ <= sub_333_2_n_31;
     end
 assign n_732 = retime_s2_22_reg_reg_IQ;
 reg retime_s2_23_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_23_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_23_reg_reg_IQ <= sub_333_2_n_55;
     end
 assign n_731 = retime_s2_23_reg_reg_IQ;
 reg retime_s2_24_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_24_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_24_reg_reg_IQ <= sub_333_2_n_59;
     end
 assign n_730 = retime_s2_24_reg_reg_IQ;
 reg retime_s2_25_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_25_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_25_reg_reg_IQ <= sub_333_2_n_7;
     end
 assign n_729 = retime_s2_25_reg_reg_IQ;
 reg retime_s2_26_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_26_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_26_reg_reg_IQ <= sub_333_2_n_8;
     end
 assign n_728 = retime_s2_26_reg_reg_IQ;
 reg retime_s2_27_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_27_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_27_reg_reg_IQ <= n_1531;
     end
 assign n_727 = retime_s2_27_reg_reg_IQ;
 reg retime_s2_28_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_28_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_28_reg_reg_IQ <= n_155;
     end
 assign n_723 = retime_s2_28_reg_reg_IQ;
 reg retime_s2_29_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_29_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_29_reg_reg_IQ <= n_101;
     end
 assign n_722 = retime_s2_29_reg_reg_IQ;
 reg retime_s2_33_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_33_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_33_reg_reg_IQ <= n_153;
     end
 assign n_716 = retime_s2_33_reg_reg_IQ;
 reg retime_s2_39_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_39_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_39_reg_reg_IQ <= n_705;
     end
 assign n_704 = retime_s2_39_reg_reg_IQ;
 reg retime_s2_40_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_40_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_40_reg_reg_IQ <= n_693;
     end
 assign n_692 = retime_s2_40_reg_reg_IQ;
 reg retime_s2_41_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_41_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_41_reg_reg_IQ <= n_683;
     end
 assign n_682 = retime_s2_41_reg_reg_IQ;
 reg retime_s2_45_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_45_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_45_reg_reg_IQ <= n_670;
     end
 assign n_669 = retime_s2_45_reg_reg_IQ;
 reg retime_s2_46_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_46_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_46_reg_reg_IQ <= n_660;
     end
 assign n_659 = retime_s2_46_reg_reg_IQ;
 reg retime_s2_48_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_48_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_48_reg_reg_IQ <= n_642;
     end
 assign n_641 = retime_s2_48_reg_reg_IQ;
 reg retime_s2_53_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_53_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_53_reg_reg_IQ <= n_628;
     end
 assign n_627 = retime_s2_53_reg_reg_IQ;
 reg retime_s2_57_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_57_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_57_reg_reg_IQ <= n_614;
     end
 assign n_613 = retime_s2_57_reg_reg_IQ;
 reg retime_s2_58_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_58_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_58_reg_reg_IQ <= n_604;
     end
 assign n_603 = retime_s2_58_reg_reg_IQ;
 reg retime_s2_59_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_59_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_59_reg_reg_IQ <= n_594;
     end
 assign n_593 = retime_s2_59_reg_reg_IQ;
 reg retime_s2_61_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_61_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_61_reg_reg_IQ <= n_192;
     end
 assign n_583 = retime_s2_61_reg_reg_IQ;
 reg retime_s2_63_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_63_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_63_reg_reg_IQ <= n_194;
     end
 assign n_581 = retime_s2_63_reg_reg_IQ;
 reg retime_s2_64_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_64_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_64_reg_reg_IQ <= n_195;
     end
 assign n_580 = retime_s2_64_reg_reg_IQ;
 reg retime_s2_65_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_65_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_65_reg_reg_IQ <= n_196;
     end
 assign n_579 = retime_s2_65_reg_reg_IQ;
 reg retime_s2_66_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_66_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_66_reg_reg_IQ <= n_197;
     end
 assign n_578 = retime_s2_66_reg_reg_IQ;
 reg retime_s2_67_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_67_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_67_reg_reg_IQ <= n_285;
     end
 assign n_577 = retime_s2_67_reg_reg_IQ;
 reg retime_s2_75_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_75_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_75_reg_reg_IQ <= n_568;
     end
 assign n_567 = retime_s2_75_reg_reg_IQ;
 reg retime_s2_76_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_76_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_76_reg_reg_IQ <= n_558;
     end
 assign n_557 = retime_s2_76_reg_reg_IQ;
 reg retime_s2_77_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_77_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_77_reg_reg_IQ <= n_548;
     end
 assign n_547 = retime_s2_77_reg_reg_IQ;
 reg retime_s2_78_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_78_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_78_reg_reg_IQ <= n_538;
     end
 assign n_537 = retime_s2_78_reg_reg_IQ;
 reg retime_s2_79_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_79_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_79_reg_reg_IQ <= n_527;
     end
 assign n_526 = retime_s2_79_reg_reg_IQ;
 reg retime_s2_90_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_90_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_90_reg_reg_IQ <= n_507;
     end
 assign n_506 = retime_s2_90_reg_reg_IQ;
 reg retime_s2_98_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_98_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_98_reg_reg_IQ <= n_486;
     end
 assign n_485 = retime_s2_98_reg_reg_IQ;
 reg retime_s2_99_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_99_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_99_reg_reg_IQ <= n_476;
     end
 assign n_475 = retime_s2_99_reg_reg_IQ;
 reg retime_s2_100_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_100_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_100_reg_reg_IQ <= n_466;
     end
 assign n_465 = retime_s2_100_reg_reg_IQ;
 reg retime_s2_101_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_101_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_101_reg_reg_IQ <= n_456;
     end
 assign n_455 = retime_s2_101_reg_reg_IQ;
 reg retime_s2_103_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_103_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_103_reg_reg_IQ <= n_445;
     end
 assign n_444 = retime_s2_103_reg_reg_IQ;
 reg retime_s2_104_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_104_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_104_reg_reg_IQ <= n_435;
     end
 assign n_434 = retime_s2_104_reg_reg_IQ;
 reg retime_s2_105_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_105_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_105_reg_reg_IQ <= n_425;
     end
 assign n_424 = retime_s2_105_reg_reg_IQ;
 reg retime_s2_106_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_106_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_106_reg_reg_IQ <= n_415;
     end
 assign n_414 = retime_s2_106_reg_reg_IQ;
 reg retime_s2_111_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_111_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_111_reg_reg_IQ <= n_401;
     end
 assign n_400 = retime_s2_111_reg_reg_IQ;
 reg retime_s2_112_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_112_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_112_reg_reg_IQ <= n_391;
     end
 assign n_390 = retime_s2_112_reg_reg_IQ;
 reg retime_s2_118_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_118_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_118_reg_reg_IQ <= n_376;
     end
 assign n_375 = retime_s2_118_reg_reg_IQ;
 reg retime_s2_120_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_120_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_120_reg_reg_IQ <= n_365;
     end
 assign n_364 = retime_s2_120_reg_reg_IQ;
 reg retime_s2_121_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_121_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_121_reg_reg_IQ <= n_355;
     end
 assign n_354 = retime_s2_121_reg_reg_IQ;
 reg retime_s2_123_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_123_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_123_reg_reg_IQ <= n_344;
     end
 assign n_343 = retime_s2_123_reg_reg_IQ;
 reg retime_s3_3_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_3_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_3_reg_reg_IQ <= n_1114;
     end
 assign n_1113 = retime_s3_3_reg_reg_IQ;
 reg retime_s3_4_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_4_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_4_reg_reg_IQ <= n_1609;
     end
 assign n_780 = retime_s3_4_reg_reg_IQ;
 reg retime_s3_5_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_5_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_5_reg_reg_IQ <= n_3257;
     end
 assign n_779 = retime_s3_5_reg_reg_IQ;
 reg retime_s3_6_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_6_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_6_reg_reg_IQ <= n_3256;
     end
 assign n_778 = retime_s3_6_reg_reg_IQ;
 reg retime_s3_7_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_7_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_7_reg_reg_IQ <= n_3258;
     end
 assign n_777 = retime_s3_7_reg_reg_IQ;
 reg retime_s3_8_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_8_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_8_reg_reg_IQ <= n_1607;
     end
 assign n_776 = retime_s3_8_reg_reg_IQ;
 reg retime_s3_9_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_9_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_9_reg_reg_IQ <= n_3049;
     end
 assign n_775 = retime_s3_9_reg_reg_IQ;
 reg retime_s3_10_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_10_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_10_reg_reg_IQ <= n_3254;
     end
 assign n_774 = retime_s3_10_reg_reg_IQ;
 reg retime_s3_11_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_11_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_11_reg_reg_IQ <= n_1601;
     end
 assign n_773 = retime_s3_11_reg_reg_IQ;
 reg retime_s3_12_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_12_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_12_reg_reg_IQ <= n_3552;
     end
 assign n_772 = retime_s3_12_reg_reg_IQ;
 reg retime_s3_13_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_13_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_13_reg_reg_IQ <= sub_390_2_n_103;
     end
 assign n_771 = retime_s3_13_reg_reg_IQ;
 reg retime_s3_14_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_14_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_14_reg_reg_IQ <= n_1614;
     end
 assign n_770 = retime_s3_14_reg_reg_IQ;
 reg retime_s3_15_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_15_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_15_reg_reg_IQ <= n_3550;
     end
 assign n_769 = retime_s3_15_reg_reg_IQ;
 reg retime_s3_16_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_16_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_16_reg_reg_IQ <= sub_390_2_n_10;
     end
 assign n_768 = retime_s3_16_reg_reg_IQ;
 reg retime_s3_17_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_17_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_17_reg_reg_IQ <= n_1599;
     end
 assign n_767 = retime_s3_17_reg_reg_IQ;
 reg retime_s3_18_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_18_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_18_reg_reg_IQ <= sub_390_2_n_59;
     end
 assign n_766 = retime_s3_18_reg_reg_IQ;
 reg retime_s3_19_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_19_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_19_reg_reg_IQ <= sub_390_2_n_36;
     end
 assign n_765 = retime_s3_19_reg_reg_IQ;
 reg retime_s3_20_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_20_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_20_reg_reg_IQ <= sub_390_2_n_19;
     end
 assign n_764 = retime_s3_20_reg_reg_IQ;
 reg retime_s3_21_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_21_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_21_reg_reg_IQ <= n_3255;
     end
 assign n_763 = retime_s3_21_reg_reg_IQ;
 reg retime_s3_22_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_22_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_22_reg_reg_IQ <= sub_390_2_n_67;
     end
 assign n_762 = retime_s3_22_reg_reg_IQ;
 reg retime_s3_23_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_23_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_23_reg_reg_IQ <= n_3261;
     end
 assign n_761 = retime_s3_23_reg_reg_IQ;
 reg retime_s3_24_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_24_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_24_reg_reg_IQ <= n_1615;
     end
 assign n_760 = retime_s3_24_reg_reg_IQ;
 reg retime_s3_25_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_25_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_25_reg_reg_IQ <= n_3259;
     end
 assign n_759 = retime_s3_25_reg_reg_IQ;
 reg retime_s3_26_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_26_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_26_reg_reg_IQ <= n_1619;
     end
 assign n_758 = retime_s3_26_reg_reg_IQ;
 reg retime_s3_27_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_27_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_27_reg_reg_IQ <= n_1616;
     end
 assign n_757 = retime_s3_27_reg_reg_IQ;
 reg retime_s3_28_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_28_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_28_reg_reg_IQ <= n_1617;
     end
 assign n_756 = retime_s3_28_reg_reg_IQ;
 reg retime_s3_29_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_29_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_29_reg_reg_IQ <= n_1618;
     end
 assign n_755 = retime_s3_29_reg_reg_IQ;
 reg retime_s3_30_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_30_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_30_reg_reg_IQ <= n_1621;
     end
 assign n_754 = retime_s3_30_reg_reg_IQ;
 reg retime_s3_31_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_31_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_31_reg_reg_IQ <= n_1620;
     end
 assign n_753 = retime_s3_31_reg_reg_IQ;
 reg retime_s3_32_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_32_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_32_reg_reg_IQ <= n_3260;
     end
 assign n_752 = retime_s3_32_reg_reg_IQ;
 reg retime_s3_33_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_33_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_33_reg_reg_IQ <= sub_390_2_n_12;
     end
 assign n_751 = retime_s3_33_reg_reg_IQ;
 reg retime_s3_36_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_36_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_36_reg_reg_IQ <= n_241;
     end
 assign n_717 = retime_s3_36_reg_reg_IQ;
 reg retime_s3_37_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_37_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_37_reg_reg_IQ <= n_242;
     end
 assign n_715 = retime_s3_37_reg_reg_IQ;
 reg retime_s3_38_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_38_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_38_reg_reg_IQ <= n_243;
     end
 assign n_714 = retime_s3_38_reg_reg_IQ;
 reg retime_s3_42_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_42_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_42_reg_reg_IQ <= n_704;
     end
 assign n_703 = retime_s3_42_reg_reg_IQ;
 reg retime_s3_43_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_43_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_43_reg_reg_IQ <= n_692;
     end
 assign n_691 = retime_s3_43_reg_reg_IQ;
 reg retime_s3_44_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_44_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_44_reg_reg_IQ <= n_682;
     end
 assign n_681 = retime_s3_44_reg_reg_IQ;
 reg retime_s3_48_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_48_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_48_reg_reg_IQ <= n_669;
     end
 assign n_668 = retime_s3_48_reg_reg_IQ;
 reg retime_s3_49_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_49_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_49_reg_reg_IQ <= n_659;
     end
 assign n_658 = retime_s3_49_reg_reg_IQ;
 reg retime_s3_51_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_51_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_51_reg_reg_IQ <= n_641;
     end
 assign n_640 = retime_s3_51_reg_reg_IQ;
 reg retime_s3_52_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_52_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_52_reg_reg_IQ <= n_252;
     end
 assign n_632 = retime_s3_52_reg_reg_IQ;
 reg retime_s3_53_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_53_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_53_reg_reg_IQ <= n_253;
     end
 assign n_631 = retime_s3_53_reg_reg_IQ;
 reg retime_s3_54_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_54_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_54_reg_reg_IQ <= n_254;
     end
 assign n_630 = retime_s3_54_reg_reg_IQ;
 reg retime_s3_56_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_56_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_56_reg_reg_IQ <= n_627;
     end
 assign n_626 = retime_s3_56_reg_reg_IQ;
 reg retime_s3_57_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_57_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_57_reg_reg_IQ <= n_256;
     end
 assign n_618 = retime_s3_57_reg_reg_IQ;
 reg retime_s3_58_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_58_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_58_reg_reg_IQ <= n_257;
     end
 assign n_616 = retime_s3_58_reg_reg_IQ;
 reg retime_s3_59_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_59_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_59_reg_reg_IQ <= n_258;
     end
 assign n_615 = retime_s3_59_reg_reg_IQ;
 reg retime_s3_60_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_60_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_60_reg_reg_IQ <= n_613;
     end
 assign n_612 = retime_s3_60_reg_reg_IQ;
 reg retime_s3_61_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_61_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_61_reg_reg_IQ <= n_603;
     end
 assign n_602 = retime_s3_61_reg_reg_IQ;
 reg retime_s3_62_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_62_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_62_reg_reg_IQ <= n_593;
     end
 assign n_592 = retime_s3_62_reg_reg_IQ;
 reg retime_s3_63_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_63_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_63_reg_reg_IQ <= n_259;
     end
 assign n_584 = retime_s3_63_reg_reg_IQ;
 reg retime_s3_64_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_64_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_64_reg_reg_IQ <= n_260;
     end
 assign n_582 = retime_s3_64_reg_reg_IQ;
 reg retime_s3_72_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_72_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_72_reg_reg_IQ <= n_567;
     end
 assign n_566 = retime_s3_72_reg_reg_IQ;
 reg retime_s3_73_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_73_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_73_reg_reg_IQ <= n_557;
     end
 assign n_556 = retime_s3_73_reg_reg_IQ;
 reg retime_s3_74_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_74_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_74_reg_reg_IQ <= n_547;
     end
 assign n_546 = retime_s3_74_reg_reg_IQ;
 reg retime_s3_75_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_75_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_75_reg_reg_IQ <= n_537;
     end
 assign n_536 = retime_s3_75_reg_reg_IQ;
 reg retime_s3_76_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_76_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_76_reg_reg_IQ <= n_526;
     end
 assign n_525 = retime_s3_76_reg_reg_IQ;
 reg retime_s3_87_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_87_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_87_reg_reg_IQ <= n_506;
     end
 assign n_505 = retime_s3_87_reg_reg_IQ;
 reg retime_s3_93_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_93_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_93_reg_reg_IQ <= n_138;
     end
 assign n_491 = retime_s3_93_reg_reg_IQ;
 reg retime_s3_95_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_95_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_95_reg_reg_IQ <= n_485;
     end
 assign n_484 = retime_s3_95_reg_reg_IQ;
 reg retime_s3_96_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_96_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_96_reg_reg_IQ <= n_475;
     end
 assign n_474 = retime_s3_96_reg_reg_IQ;
 reg retime_s3_97_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_97_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_97_reg_reg_IQ <= n_465;
     end
 assign n_464 = retime_s3_97_reg_reg_IQ;
 reg retime_s3_98_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_98_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_98_reg_reg_IQ <= n_455;
     end
 assign n_454 = retime_s3_98_reg_reg_IQ;
 reg retime_s3_100_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_100_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_100_reg_reg_IQ <= n_444;
     end
 assign n_443 = retime_s3_100_reg_reg_IQ;
 reg retime_s3_101_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_101_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_101_reg_reg_IQ <= n_434;
     end
 assign n_433 = retime_s3_101_reg_reg_IQ;
 reg retime_s3_102_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_102_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_102_reg_reg_IQ <= n_424;
     end
 assign n_423 = retime_s3_102_reg_reg_IQ;
 reg retime_s3_103_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_103_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_103_reg_reg_IQ <= n_414;
     end
 assign n_413 = retime_s3_103_reg_reg_IQ;
 reg retime_s3_108_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_108_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_108_reg_reg_IQ <= n_400;
     end
 assign n_399 = retime_s3_108_reg_reg_IQ;
 reg retime_s3_109_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_109_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_109_reg_reg_IQ <= n_390;
     end
 assign n_389 = retime_s3_109_reg_reg_IQ;
 reg retime_s3_115_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_115_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_115_reg_reg_IQ <= n_375;
     end
 assign n_374 = retime_s3_115_reg_reg_IQ;
 reg retime_s3_117_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_117_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_117_reg_reg_IQ <= n_364;
     end
 assign n_363 = retime_s3_117_reg_reg_IQ;
 reg retime_s3_118_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_118_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_118_reg_reg_IQ <= n_354;
     end
 assign n_353 = retime_s3_118_reg_reg_IQ;
 reg retime_s3_120_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_120_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_120_reg_reg_IQ <= n_343;
     end
 assign n_342 = retime_s3_120_reg_reg_IQ;
 reg retime_s4_3_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_3_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_3_reg_reg_IQ <= n_1113;
     end
 assign n_1112 = retime_s4_3_reg_reg_IQ;
 reg retime_s4_4_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_4_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_4_reg_reg_IQ <= n_3295;
     end
 assign n_832 = retime_s4_4_reg_reg_IQ;
 reg retime_s4_5_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_5_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_5_reg_reg_IQ <= sub_466_2_n_87;
     end
 assign n_831 = retime_s4_5_reg_reg_IQ;
 reg retime_s4_6_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_6_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_6_reg_reg_IQ <= sub_466_2_n_84;
     end
 assign n_830 = retime_s4_6_reg_reg_IQ;
 reg retime_s4_7_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_7_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_7_reg_reg_IQ <= sub_466_2_n_15;
     end
 assign n_829 = retime_s4_7_reg_reg_IQ;
 reg retime_s4_8_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_8_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_8_reg_reg_IQ <= n_3299;
     end
 assign n_828 = retime_s4_8_reg_reg_IQ;
 reg retime_s4_9_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_9_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_9_reg_reg_IQ <= n_3306;
     end
 assign n_827 = retime_s4_9_reg_reg_IQ;
 reg retime_s4_10_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_10_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_10_reg_reg_IQ <= sub_466_2_n_39;
     end
 assign n_826 = retime_s4_10_reg_reg_IQ;
 reg retime_s4_11_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_11_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_11_reg_reg_IQ <= sub_466_2_n_58;
     end
 assign n_825 = retime_s4_11_reg_reg_IQ;
 reg retime_s4_12_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_12_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_12_reg_reg_IQ <= sub_466_2_n_14;
     end
 assign n_824 = retime_s4_12_reg_reg_IQ;
 reg retime_s4_13_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_13_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_13_reg_reg_IQ <= sub_466_2_n_74;
     end
 assign n_823 = retime_s4_13_reg_reg_IQ;
 reg retime_s4_14_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_14_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_14_reg_reg_IQ <= sub_466_2_n_88;
     end
 assign n_822 = retime_s4_14_reg_reg_IQ;
 reg retime_s4_15_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_15_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_15_reg_reg_IQ <= n_3294;
     end
 assign n_821 = retime_s4_15_reg_reg_IQ;
 reg retime_s4_16_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_16_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_16_reg_reg_IQ <= n_3296;
     end
 assign n_820 = retime_s4_16_reg_reg_IQ;
 reg retime_s4_17_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_17_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_17_reg_reg_IQ <= sub_466_2_n_9;
     end
 assign n_819 = retime_s4_17_reg_reg_IQ;
 reg retime_s4_18_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_18_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_18_reg_reg_IQ <= sub_466_2_n_89;
     end
 assign n_818 = retime_s4_18_reg_reg_IQ;
 reg retime_s4_19_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_19_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_19_reg_reg_IQ <= sub_466_2_n_17;
     end
 assign n_817 = retime_s4_19_reg_reg_IQ;
 reg retime_s4_20_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_20_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_20_reg_reg_IQ <= sub_466_2_n_46;
     end
 assign n_816 = retime_s4_20_reg_reg_IQ;
 reg retime_s4_21_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_21_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_21_reg_reg_IQ <= sub_466_2_n_85;
     end
 assign n_815 = retime_s4_21_reg_reg_IQ;
 reg retime_s4_22_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_22_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_22_reg_reg_IQ <= sub_466_2_n_12;
     end
 assign n_814 = retime_s4_22_reg_reg_IQ;
 reg retime_s4_23_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_23_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_23_reg_reg_IQ <= sub_466_2_n_71;
     end
 assign n_813 = retime_s4_23_reg_reg_IQ;
 reg retime_s4_24_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_24_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_24_reg_reg_IQ <= n_3297;
     end
 assign n_812 = retime_s4_24_reg_reg_IQ;
 reg retime_s4_25_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_25_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_25_reg_reg_IQ <= sub_466_2_n_10;
     end
 assign n_811 = retime_s4_25_reg_reg_IQ;
 reg retime_s4_26_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_26_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_26_reg_reg_IQ <= sub_466_2_n_65;
     end
 assign n_810 = retime_s4_26_reg_reg_IQ;
 reg retime_s4_27_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_27_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_27_reg_reg_IQ <= n_1725;
     end
 assign n_809 = retime_s4_27_reg_reg_IQ;
 reg retime_s4_28_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_28_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_28_reg_reg_IQ <= sub_466_2_n_1;
     end
 assign n_808 = retime_s4_28_reg_reg_IQ;
 reg retime_s4_29_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_29_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_29_reg_reg_IQ <= sub_466_2_n_25;
     end
 assign n_807 = retime_s4_29_reg_reg_IQ;
 reg retime_s4_30_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_30_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_30_reg_reg_IQ <= n_3298;
     end
 assign n_806 = retime_s4_30_reg_reg_IQ;
 reg retime_s4_31_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_31_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_31_reg_reg_IQ <= n_3301;
     end
 assign n_805 = retime_s4_31_reg_reg_IQ;
 reg retime_s4_32_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_32_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_32_reg_reg_IQ <= sub_466_2_n_7;
     end
 assign n_804 = retime_s4_32_reg_reg_IQ;
 reg retime_s4_33_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_33_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_33_reg_reg_IQ <= sub_466_2_n_79;
     end
 assign n_803 = retime_s4_33_reg_reg_IQ;
 reg retime_s4_34_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_34_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_34_reg_reg_IQ <= sub_466_2_n_67;
     end
 assign n_802 = retime_s4_34_reg_reg_IQ;
 reg retime_s4_35_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_35_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_35_reg_reg_IQ <= sub_466_2_n_86;
     end
 assign n_801 = retime_s4_35_reg_reg_IQ;
 reg retime_s4_36_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_36_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_36_reg_reg_IQ <= n_3302;
     end
 assign n_800 = retime_s4_36_reg_reg_IQ;
 reg retime_s4_37_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_37_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_37_reg_reg_IQ <= n_3303;
     end
 assign n_799 = retime_s4_37_reg_reg_IQ;
 reg retime_s4_38_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_38_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_38_reg_reg_IQ <= sub_466_2_n_73;
     end
 assign n_798 = retime_s4_38_reg_reg_IQ;
 reg retime_s4_39_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_39_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_39_reg_reg_IQ <= sub_466_2_n_6;
     end
 assign n_797 = retime_s4_39_reg_reg_IQ;
 reg retime_s4_40_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_40_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_40_reg_reg_IQ <= sub_466_2_n_44;
     end
 assign n_796 = retime_s4_40_reg_reg_IQ;
 reg retime_s4_41_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_41_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_41_reg_reg_IQ <= n_3304;
     end
 assign n_795 = retime_s4_41_reg_reg_IQ;
 reg retime_s4_42_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_42_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_42_reg_reg_IQ <= n_3305;
     end
 assign n_794 = retime_s4_42_reg_reg_IQ;
 reg retime_s4_43_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_43_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_43_reg_reg_IQ <= sub_466_2_n_8;
     end
 assign n_793 = retime_s4_43_reg_reg_IQ;
 reg retime_s4_44_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_44_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_44_reg_reg_IQ <= sub_466_2_n_41;
     end
 assign n_792 = retime_s4_44_reg_reg_IQ;
 reg retime_s4_45_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_45_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_45_reg_reg_IQ <= sub_466_2_n_0;
     end
 assign n_791 = retime_s4_45_reg_reg_IQ;
 reg retime_s4_46_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_46_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_46_reg_reg_IQ <= sub_466_2_n_55;
     end
 assign n_790 = retime_s4_46_reg_reg_IQ;
 reg retime_s4_47_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_47_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_47_reg_reg_IQ <= n_1727;
     end
 assign n_789 = retime_s4_47_reg_reg_IQ;
 reg retime_s4_48_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_48_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_48_reg_reg_IQ <= sub_466_2_n_102;
     end
 assign n_788 = retime_s4_48_reg_reg_IQ;
 reg retime_s4_49_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_49_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_49_reg_reg_IQ <= n_1744;
     end
 assign n_787 = retime_s4_49_reg_reg_IQ;
 reg retime_s4_50_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_50_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_50_reg_reg_IQ <= n_1728;
     end
 assign n_786 = retime_s4_50_reg_reg_IQ;
 reg retime_s4_51_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_51_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_51_reg_reg_IQ <= n_1745;
     end
 assign n_785 = retime_s4_51_reg_reg_IQ;
 reg retime_s4_52_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_52_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_52_reg_reg_IQ <= sub_466_2_n_49;
     end
 assign n_784 = retime_s4_52_reg_reg_IQ;
 reg retime_s4_53_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_53_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_53_reg_reg_IQ <= n_3300;
     end
 assign n_783 = retime_s4_53_reg_reg_IQ;
 reg retime_s4_54_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_54_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_54_reg_reg_IQ <= sub_466_2_n_76;
     end
 assign n_782 = retime_s4_54_reg_reg_IQ;
 reg retime_s4_55_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_55_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_55_reg_reg_IQ <= sub_466_2_n_105;
     end
 assign n_781 = retime_s4_55_reg_reg_IQ;
 reg retime_s4_56_reg_reg_IQ;
 wire retime_s4_56_reg_reg_IQN;
 assign retime_s4_56_reg_reg_IQN = !retime_s4_56_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_56_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_56_reg_reg_IQ <= n_24;
     end
 assign n_299 = retime_s4_56_reg_reg_IQN;
 reg retime_s4_57_reg_reg_IQ;
 wire retime_s4_57_reg_reg_IQN;
 assign retime_s4_57_reg_reg_IQN = !retime_s4_57_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_57_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_57_reg_reg_IQ <= n_171;
     end
 assign n_297 = retime_s4_57_reg_reg_IQN;
 reg retime_s4_58_reg_reg_IQ;
 wire retime_s4_58_reg_reg_IQN;
 assign retime_s4_58_reg_reg_IQN = !retime_s4_58_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_58_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_58_reg_reg_IQ <= n_23;
     end
 assign n_295 = retime_s4_58_reg_reg_IQN;
 reg retime_s4_59_reg_reg_IQ;
 wire retime_s4_59_reg_reg_IQN;
 assign retime_s4_59_reg_reg_IQN = !retime_s4_59_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_59_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_59_reg_reg_IQ <= n_174;
     end
 assign n_293 = retime_s4_59_reg_reg_IQN;
 reg retime_s4_61_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_61_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_61_reg_reg_IQ <= n_703;
     end
 assign n_702 = retime_s4_61_reg_reg_IQ;
 reg retime_s4_62_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_62_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_62_reg_reg_IQ <= n_691;
     end
 assign n_690 = retime_s4_62_reg_reg_IQ;
 reg retime_s4_63_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_63_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_63_reg_reg_IQ <= n_681;
     end
 assign n_680 = retime_s4_63_reg_reg_IQ;
 reg retime_s4_64_reg_reg_IQ;
 wire retime_s4_64_reg_reg_IQN;
 assign retime_s4_64_reg_reg_IQN = !retime_s4_64_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_64_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_64_reg_reg_IQ <= n_67;
     end
 assign n_289 = retime_s4_64_reg_reg_IQN;
 reg retime_s4_66_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_66_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_66_reg_reg_IQ <= n_66;
     end
 assign n_671 = retime_s4_66_reg_reg_IQ;
 reg retime_s4_67_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_67_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_67_reg_reg_IQ <= n_668;
     end
 assign n_667 = retime_s4_67_reg_reg_IQ;
 reg retime_s4_68_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_68_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_68_reg_reg_IQ <= n_658;
     end
 assign n_657 = retime_s4_68_reg_reg_IQ;
 reg retime_s4_69_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_69_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_69_reg_reg_IQ <= n_124;
     end
 assign n_650 = retime_s4_69_reg_reg_IQ;
 reg retime_s4_70_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_70_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_70_reg_reg_IQ <= n_640;
     end
 assign n_639 = retime_s4_70_reg_reg_IQ;
 reg retime_s4_71_reg_reg_IQ;
 wire retime_s4_71_reg_reg_IQN;
 assign retime_s4_71_reg_reg_IQN = !retime_s4_71_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_71_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_71_reg_reg_IQ <= n_22;
     end
 assign n_286 = retime_s4_71_reg_reg_IQN;
 reg retime_s4_72_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_72_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_72_reg_reg_IQ <= n_626;
     end
 assign n_625 = retime_s4_72_reg_reg_IQ;
 reg retime_s4_73_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_73_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_73_reg_reg_IQ <= n_612;
     end
 assign n_611 = retime_s4_73_reg_reg_IQ;
 reg retime_s4_74_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_74_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_74_reg_reg_IQ <= n_602;
     end
 assign n_601 = retime_s4_74_reg_reg_IQ;
 reg retime_s4_75_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_75_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_75_reg_reg_IQ <= n_592;
     end
 assign n_591 = retime_s4_75_reg_reg_IQ;
 reg retime_s4_83_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_83_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_83_reg_reg_IQ <= n_566;
     end
 assign n_565 = retime_s4_83_reg_reg_IQ;
 reg retime_s4_84_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_84_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_84_reg_reg_IQ <= n_556;
     end
 assign n_555 = retime_s4_84_reg_reg_IQ;
 reg retime_s4_85_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_85_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_85_reg_reg_IQ <= n_546;
     end
 assign n_545 = retime_s4_85_reg_reg_IQ;
 reg retime_s4_86_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_86_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_86_reg_reg_IQ <= n_536;
     end
 assign n_535 = retime_s4_86_reg_reg_IQ;
 reg retime_s4_87_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_87_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_87_reg_reg_IQ <= n_525;
     end
 assign n_524 = retime_s4_87_reg_reg_IQ;
 reg retime_s4_98_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_98_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_98_reg_reg_IQ <= n_505;
     end
 assign n_504 = retime_s4_98_reg_reg_IQ;
 reg retime_s4_103_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_103_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_103_reg_reg_IQ <= n_116;
     end
 assign n_492 = retime_s4_103_reg_reg_IQ;
 reg retime_s4_104_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_104_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_104_reg_reg_IQ <= n_55;
     end
 assign n_490 = retime_s4_104_reg_reg_IQ;
 reg retime_s4_105_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_105_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_105_reg_reg_IQ <= n_484;
     end
 assign n_483 = retime_s4_105_reg_reg_IQ;
 reg retime_s4_106_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_106_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_106_reg_reg_IQ <= n_474;
     end
 assign n_473 = retime_s4_106_reg_reg_IQ;
 reg retime_s4_107_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_107_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_107_reg_reg_IQ <= n_464;
     end
 assign n_463 = retime_s4_107_reg_reg_IQ;
 reg retime_s4_108_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_108_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_108_reg_reg_IQ <= n_454;
     end
 assign n_453 = retime_s4_108_reg_reg_IQ;
 reg retime_s4_110_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_110_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_110_reg_reg_IQ <= n_443;
     end
 assign n_442 = retime_s4_110_reg_reg_IQ;
 reg retime_s4_111_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_111_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_111_reg_reg_IQ <= n_433;
     end
 assign n_432 = retime_s4_111_reg_reg_IQ;
 reg retime_s4_112_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_112_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_112_reg_reg_IQ <= n_423;
     end
 assign n_422 = retime_s4_112_reg_reg_IQ;
 reg retime_s4_113_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_113_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_113_reg_reg_IQ <= n_413;
     end
 assign n_412 = retime_s4_113_reg_reg_IQ;
 reg retime_s4_114_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_114_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_114_reg_reg_IQ <= n_52;
     end
 assign n_405 = retime_s4_114_reg_reg_IQ;
 reg retime_s4_115_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_115_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_115_reg_reg_IQ <= n_53;
     end
 assign n_404 = retime_s4_115_reg_reg_IQ;
 reg retime_s4_116_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_116_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_116_reg_reg_IQ <= n_54;
     end
 assign n_403 = retime_s4_116_reg_reg_IQ;
 reg retime_s4_117_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_117_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_117_reg_reg_IQ <= n_127;
     end
 assign n_402 = retime_s4_117_reg_reg_IQ;
 reg retime_s4_118_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_118_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_118_reg_reg_IQ <= n_399;
     end
 assign n_398 = retime_s4_118_reg_reg_IQ;
 reg retime_s4_119_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_119_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_119_reg_reg_IQ <= n_389;
     end
 assign n_388 = retime_s4_119_reg_reg_IQ;
 reg retime_s4_120_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_120_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_120_reg_reg_IQ <= n_50;
     end
 assign n_381 = retime_s4_120_reg_reg_IQ;
 reg retime_s4_125_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_125_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_125_reg_reg_IQ <= n_374;
     end
 assign n_373 = retime_s4_125_reg_reg_IQ;
 reg retime_s4_127_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_127_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_127_reg_reg_IQ <= n_363;
     end
 assign n_362 = retime_s4_127_reg_reg_IQ;
 reg retime_s4_128_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_128_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_128_reg_reg_IQ <= n_353;
     end
 assign n_352 = retime_s4_128_reg_reg_IQ;
 reg retime_s4_130_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_130_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_130_reg_reg_IQ <= n_342;
     end
 assign n_341 = retime_s4_130_reg_reg_IQ;
 reg retime_s5_3_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_3_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_3_reg_reg_IQ <= n_1112;
     end
 assign n_1111 = retime_s5_3_reg_reg_IQ;
 reg retime_s5_4_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_4_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_4_reg_reg_IQ <= n_3338;
     end
 assign n_853 = retime_s5_4_reg_reg_IQ;
 reg retime_s5_5_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_5_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_5_reg_reg_IQ <= n_3331;
     end
 assign n_852 = retime_s5_5_reg_reg_IQ;
 reg retime_s5_6_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_6_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_6_reg_reg_IQ <= n_3337;
     end
 assign n_851 = retime_s5_6_reg_reg_IQ;
 reg retime_s5_7_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_7_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_7_reg_reg_IQ <= n_3332;
     end
 assign n_850 = retime_s5_7_reg_reg_IQ;
 reg retime_s5_8_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_8_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_8_reg_reg_IQ <= n_3333;
     end
 assign n_849 = retime_s5_8_reg_reg_IQ;
 reg retime_s5_9_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_9_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_9_reg_reg_IQ <= n_3339;
     end
 assign n_848 = retime_s5_9_reg_reg_IQ;
 reg retime_s5_10_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_10_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_10_reg_reg_IQ <= n_3341;
     end
 assign n_847 = retime_s5_10_reg_reg_IQ;
 reg retime_s5_11_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_11_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_11_reg_reg_IQ <= n_3736;
     end
 assign n_846 = retime_s5_11_reg_reg_IQ;
 reg retime_s5_12_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_12_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_12_reg_reg_IQ <= n_3738;
     end
 assign n_845 = retime_s5_12_reg_reg_IQ;
 reg retime_s5_13_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_13_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_13_reg_reg_IQ <= n_3744;
     end
 assign n_844 = retime_s5_13_reg_reg_IQ;
 reg retime_s5_14_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_14_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_14_reg_reg_IQ <= n_3059;
     end
 assign n_843 = retime_s5_14_reg_reg_IQ;
 reg retime_s5_15_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_15_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_15_reg_reg_IQ <= n_3741;
     end
 assign n_842 = retime_s5_15_reg_reg_IQ;
 reg retime_s5_16_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_16_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_16_reg_reg_IQ <= n_3740;
     end
 assign n_841 = retime_s5_16_reg_reg_IQ;
 reg retime_s5_17_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_17_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_17_reg_reg_IQ <= sub_523_2_n_107;
     end
 assign n_840 = retime_s5_17_reg_reg_IQ;
 reg retime_s5_18_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_18_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_18_reg_reg_IQ <= n_1859;
     end
 assign n_839 = retime_s5_18_reg_reg_IQ;
 reg retime_s5_19_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_19_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_19_reg_reg_IQ <= n_3739;
     end
 assign n_838 = retime_s5_19_reg_reg_IQ;
 reg retime_s5_20_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_20_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_20_reg_reg_IQ <= n_3743;
     end
 assign n_837 = retime_s5_20_reg_reg_IQ;
 reg retime_s5_21_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_21_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_21_reg_reg_IQ <= n_3737;
     end
 assign n_836 = retime_s5_21_reg_reg_IQ;
 reg retime_s5_22_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_22_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_22_reg_reg_IQ <= n_1828;
     end
 assign n_835 = retime_s5_22_reg_reg_IQ;
 reg retime_s5_23_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_23_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_23_reg_reg_IQ <= n_3742;
     end
 assign n_834 = retime_s5_23_reg_reg_IQ;
 reg retime_s5_24_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_24_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_24_reg_reg_IQ <= n_3735;
     end
 assign n_833 = retime_s5_24_reg_reg_IQ;
 reg retime_s5_25_reg_reg_IQ;
 wire retime_s5_25_reg_reg_IQN;
 assign retime_s5_25_reg_reg_IQN = !retime_s5_25_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_25_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_25_reg_reg_IQ <= n_299;
     end
 assign n_298 = retime_s5_25_reg_reg_IQN;
 reg retime_s5_26_reg_reg_IQ;
 wire retime_s5_26_reg_reg_IQN;
 assign retime_s5_26_reg_reg_IQN = !retime_s5_26_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_26_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_26_reg_reg_IQ <= n_297;
     end
 assign n_296 = retime_s5_26_reg_reg_IQN;
 reg retime_s5_27_reg_reg_IQ;
 wire retime_s5_27_reg_reg_IQN;
 assign retime_s5_27_reg_reg_IQN = !retime_s5_27_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_27_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_27_reg_reg_IQ <= n_295;
     end
 assign n_294 = retime_s5_27_reg_reg_IQN;
 reg retime_s5_28_reg_reg_IQ;
 wire retime_s5_28_reg_reg_IQN;
 assign retime_s5_28_reg_reg_IQN = !retime_s5_28_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_28_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_28_reg_reg_IQ <= n_293;
     end
 assign n_709 = retime_s5_28_reg_reg_IQN;
 reg retime_s5_29_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_29_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_29_reg_reg_IQ <= n_9;
     end
 assign n_292 = retime_s5_29_reg_reg_IQ;
 reg retime_s5_30_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_30_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_30_reg_reg_IQ <= n_702;
     end
 assign n_701 = retime_s5_30_reg_reg_IQ;
 reg retime_s5_31_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_31_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_31_reg_reg_IQ <= n_690;
     end
 assign n_689 = retime_s5_31_reg_reg_IQ;
 reg retime_s5_32_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_32_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_32_reg_reg_IQ <= n_680;
     end
 assign n_679 = retime_s5_32_reg_reg_IQ;
 reg retime_s5_33_reg_reg_IQ;
 wire retime_s5_33_reg_reg_IQN;
 assign retime_s5_33_reg_reg_IQN = !retime_s5_33_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_33_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_33_reg_reg_IQ <= n_289;
     end
 assign n_288 = retime_s5_33_reg_reg_IQN;
 reg retime_s5_34_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_34_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_34_reg_reg_IQ <= n_119;
     end
 assign n_287 = retime_s5_34_reg_reg_IQ;
 reg retime_s5_35_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_35_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_35_reg_reg_IQ <= n_667;
     end
 assign n_666 = retime_s5_35_reg_reg_IQ;
 reg retime_s5_36_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_36_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_36_reg_reg_IQ <= n_657;
     end
 assign n_656 = retime_s5_36_reg_reg_IQ;
 reg retime_s5_37_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_37_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_37_reg_reg_IQ <= n_639;
     end
 assign n_638 = retime_s5_37_reg_reg_IQ;
 reg retime_s5_38_reg_reg_IQ;
 wire retime_s5_38_reg_reg_IQN;
 assign retime_s5_38_reg_reg_IQN = !retime_s5_38_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_38_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_38_reg_reg_IQ <= n_286;
     end
 assign n_629 = retime_s5_38_reg_reg_IQN;
 reg retime_s5_39_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_39_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_39_reg_reg_IQ <= n_625;
     end
 assign n_624 = retime_s5_39_reg_reg_IQ;
 reg retime_s5_40_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_40_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_40_reg_reg_IQ <= n_611;
     end
 assign n_610 = retime_s5_40_reg_reg_IQ;
 reg retime_s5_41_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_41_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_41_reg_reg_IQ <= n_601;
     end
 assign n_600 = retime_s5_41_reg_reg_IQ;
 reg retime_s5_42_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_42_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_42_reg_reg_IQ <= n_591;
     end
 assign n_590 = retime_s5_42_reg_reg_IQ;
 reg retime_s5_43_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_43_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_43_reg_reg_IQ <= n_45;
     end
 assign n_575 = retime_s5_43_reg_reg_IQ;
 reg retime_s5_48_reg_reg_IQ;
 wire retime_s5_48_reg_reg_IQN;
 assign retime_s5_48_reg_reg_IQN = !retime_s5_48_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_48_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_48_reg_reg_IQ <= n_165;
     end
 assign n_284 = retime_s5_48_reg_reg_IQN;
 reg retime_s5_49_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_49_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_49_reg_reg_IQ <= n_164;
     end
 assign n_281 = retime_s5_49_reg_reg_IQ;
 reg retime_s5_50_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_50_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_50_reg_reg_IQ <= n_565;
     end
 assign n_564 = retime_s5_50_reg_reg_IQ;
 reg retime_s5_51_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_51_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_51_reg_reg_IQ <= n_555;
     end
 assign n_554 = retime_s5_51_reg_reg_IQ;
 reg retime_s5_52_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_52_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_52_reg_reg_IQ <= n_545;
     end
 assign n_544 = retime_s5_52_reg_reg_IQ;
 reg retime_s5_53_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_53_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_53_reg_reg_IQ <= n_535;
     end
 assign n_534 = retime_s5_53_reg_reg_IQ;
 reg retime_s5_54_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_54_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_54_reg_reg_IQ <= n_524;
     end
 assign n_523 = retime_s5_54_reg_reg_IQ;
 reg retime_s5_57_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_57_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_57_reg_reg_IQ <= n_120;
     end
 assign n_280 = retime_s5_57_reg_reg_IQ;
 reg retime_s5_60_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_60_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_60_reg_reg_IQ <= n_43;
     end
 assign n_278 = retime_s5_60_reg_reg_IQ;
 reg retime_s5_64_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_64_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_64_reg_reg_IQ <= n_41;
     end
 assign n_277 = retime_s5_64_reg_reg_IQ;
 reg retime_s5_65_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_65_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_65_reg_reg_IQ <= n_504;
     end
 assign n_503 = retime_s5_65_reg_reg_IQ;
 reg retime_s5_67_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_67_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_67_reg_reg_IQ <= n_108;
     end
 assign n_496 = retime_s5_67_reg_reg_IQ;
 reg retime_s5_68_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_68_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_68_reg_reg_IQ <= n_6;
     end
 assign n_495 = retime_s5_68_reg_reg_IQ;
 reg retime_s5_69_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_69_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_69_reg_reg_IQ <= n_73;
     end
 assign n_493 = retime_s5_69_reg_reg_IQ;
 reg retime_s5_70_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_70_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_70_reg_reg_IQ <= n_483;
     end
 assign n_482 = retime_s5_70_reg_reg_IQ;
 reg retime_s5_71_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_71_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_71_reg_reg_IQ <= n_473;
     end
 assign n_472 = retime_s5_71_reg_reg_IQ;
 reg retime_s5_72_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_72_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_72_reg_reg_IQ <= n_463;
     end
 assign n_462 = retime_s5_72_reg_reg_IQ;
 reg retime_s5_73_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_73_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_73_reg_reg_IQ <= n_453;
     end
 assign n_452 = retime_s5_73_reg_reg_IQ;
 reg retime_s5_74_reg_reg_IQ;
 wire retime_s5_74_reg_reg_IQN;
 assign retime_s5_74_reg_reg_IQN = !retime_s5_74_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_74_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_74_reg_reg_IQ <= n_5;
     end
 assign n_273 = retime_s5_74_reg_reg_IQN;
 reg retime_s5_75_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_75_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_75_reg_reg_IQ <= n_442;
     end
 assign n_441 = retime_s5_75_reg_reg_IQ;
 reg retime_s5_76_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_76_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_76_reg_reg_IQ <= n_432;
     end
 assign n_431 = retime_s5_76_reg_reg_IQ;
 reg retime_s5_77_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_77_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_77_reg_reg_IQ <= n_422;
     end
 assign n_421 = retime_s5_77_reg_reg_IQ;
 reg retime_s5_78_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_78_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_78_reg_reg_IQ <= n_412;
     end
 assign n_411 = retime_s5_78_reg_reg_IQ;
 reg retime_s5_79_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_79_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_79_reg_reg_IQ <= n_398;
     end
 assign n_397 = retime_s5_79_reg_reg_IQ;
 reg retime_s5_80_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_80_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_80_reg_reg_IQ <= n_388;
     end
 assign n_387 = retime_s5_80_reg_reg_IQ;
 reg retime_s5_82_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_82_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_82_reg_reg_IQ <= n_158;
     end
 assign n_271 = retime_s5_82_reg_reg_IQ;
 reg retime_s5_84_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_84_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_84_reg_reg_IQ <= n_157;
     end
 assign n_269 = retime_s5_84_reg_reg_IQ;
 reg retime_s5_85_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_85_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_85_reg_reg_IQ <= n_373;
     end
 assign n_372 = retime_s5_85_reg_reg_IQ;
 reg retime_s5_87_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_87_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_87_reg_reg_IQ <= n_362;
     end
 assign n_361 = retime_s5_87_reg_reg_IQ;
 reg retime_s5_88_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_88_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_88_reg_reg_IQ <= n_352;
     end
 assign n_351 = retime_s5_88_reg_reg_IQ;
 reg retime_s5_90_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_90_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_90_reg_reg_IQ <= n_341;
     end
 assign n_340 = retime_s5_90_reg_reg_IQ;
 reg retime_s6_3_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_3_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_3_reg_reg_IQ <= n_1111;
     end
 assign n_1110 = retime_s6_3_reg_reg_IQ;
 reg retime_s6_4_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_4_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_4_reg_reg_IQ <= n_3363;
     end
 assign n_912 = retime_s6_4_reg_reg_IQ;
 reg retime_s6_5_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_5_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_5_reg_reg_IQ <= n_3366;
     end
 assign n_911 = retime_s6_5_reg_reg_IQ;
 reg retime_s6_6_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_6_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_6_reg_reg_IQ <= sub_561_2_n_67;
     end
 assign n_910 = retime_s6_6_reg_reg_IQ;
 reg retime_s6_7_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_7_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_7_reg_reg_IQ <= n_3365;
     end
 assign n_909 = retime_s6_7_reg_reg_IQ;
 reg retime_s6_8_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_8_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_8_reg_reg_IQ <= sub_561_2_n_17;
     end
 assign n_908 = retime_s6_8_reg_reg_IQ;
 reg retime_s6_9_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_9_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_9_reg_reg_IQ <= sub_561_2_n_66;
     end
 assign n_907 = retime_s6_9_reg_reg_IQ;
 reg retime_s6_10_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_10_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_10_reg_reg_IQ <= n_3614;
     end
 assign n_906 = retime_s6_10_reg_reg_IQ;
 reg retime_s6_11_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_11_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_11_reg_reg_IQ <= sub_561_2_n_16;
     end
 assign n_905 = retime_s6_11_reg_reg_IQ;
 reg retime_s6_12_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_12_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_12_reg_reg_IQ <= sub_561_2_n_122;
     end
 assign n_904 = retime_s6_12_reg_reg_IQ;
 reg retime_s6_13_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_13_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_13_reg_reg_IQ <= sub_561_2_n_110;
     end
 assign n_903 = retime_s6_13_reg_reg_IQ;
 reg retime_s6_14_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_14_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_14_reg_reg_IQ <= n_3375;
     end
 assign n_902 = retime_s6_14_reg_reg_IQ;
 reg retime_s6_15_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_15_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_15_reg_reg_IQ <= n_3380;
     end
 assign n_901 = retime_s6_15_reg_reg_IQ;
 reg retime_s6_16_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_16_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_16_reg_reg_IQ <= n_3373;
     end
 assign n_900 = retime_s6_16_reg_reg_IQ;
 reg retime_s6_17_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_17_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_17_reg_reg_IQ <= sub_561_2_n_4;
     end
 assign n_899 = retime_s6_17_reg_reg_IQ;
 reg retime_s6_18_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_18_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_18_reg_reg_IQ <= sub_561_2_n_152;
     end
 assign n_898 = retime_s6_18_reg_reg_IQ;
 reg retime_s6_19_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_19_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_19_reg_reg_IQ <= sub_561_2_n_106;
     end
 assign n_897 = retime_s6_19_reg_reg_IQ;
 reg retime_s6_20_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_20_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_20_reg_reg_IQ <= n_1936;
     end
 assign n_896 = retime_s6_20_reg_reg_IQ;
 reg retime_s6_21_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_21_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_21_reg_reg_IQ <= sub_561_2_n_65;
     end
 assign n_895 = retime_s6_21_reg_reg_IQ;
 reg retime_s6_22_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_22_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_22_reg_reg_IQ <= n_3615;
     end
 assign n_894 = retime_s6_22_reg_reg_IQ;
 reg retime_s6_23_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_23_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_23_reg_reg_IQ <= sub_561_2_n_112;
     end
 assign n_893 = retime_s6_23_reg_reg_IQ;
 reg retime_s6_24_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_24_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_24_reg_reg_IQ <= sub_561_2_n_96;
     end
 assign n_892 = retime_s6_24_reg_reg_IQ;
 reg retime_s6_25_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_25_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_25_reg_reg_IQ <= n_3618;
     end
 assign n_891 = retime_s6_25_reg_reg_IQ;
 reg retime_s6_26_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_26_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_26_reg_reg_IQ <= sub_561_2_n_92;
     end
 assign n_890 = retime_s6_26_reg_reg_IQ;
 reg retime_s6_27_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_27_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_27_reg_reg_IQ <= n_1916;
     end
 assign n_889 = retime_s6_27_reg_reg_IQ;
 reg retime_s6_28_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_28_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_28_reg_reg_IQ <= n_3364;
     end
 assign n_888 = retime_s6_28_reg_reg_IQ;
 reg retime_s6_29_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_29_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_29_reg_reg_IQ <= sub_561_2_n_63;
     end
 assign n_887 = retime_s6_29_reg_reg_IQ;
 reg retime_s6_30_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_30_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_30_reg_reg_IQ <= sub_561_2_n_24;
     end
 assign n_886 = retime_s6_30_reg_reg_IQ;
 reg retime_s6_31_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_31_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_31_reg_reg_IQ <= sub_561_2_n_58;
     end
 assign n_885 = retime_s6_31_reg_reg_IQ;
 reg retime_s6_32_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_32_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_32_reg_reg_IQ <= n_1938;
     end
 assign n_884 = retime_s6_32_reg_reg_IQ;
 reg retime_s6_33_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_33_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_33_reg_reg_IQ <= n_1937;
     end
 assign n_883 = retime_s6_33_reg_reg_IQ;
 reg retime_s6_34_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_34_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_34_reg_reg_IQ <= n_3367;
     end
 assign n_882 = retime_s6_34_reg_reg_IQ;
 reg retime_s6_35_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_35_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_35_reg_reg_IQ <= n_3368;
     end
 assign n_881 = retime_s6_35_reg_reg_IQ;
 reg retime_s6_36_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_36_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_36_reg_reg_IQ <= n_1939;
     end
 assign n_880 = retime_s6_36_reg_reg_IQ;
 reg retime_s6_37_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_37_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_37_reg_reg_IQ <= n_1940;
     end
 assign n_879 = retime_s6_37_reg_reg_IQ;
 reg retime_s6_38_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_38_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_38_reg_reg_IQ <= n_3369;
     end
 assign n_878 = retime_s6_38_reg_reg_IQ;
 reg retime_s6_39_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_39_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_39_reg_reg_IQ <= n_3370;
     end
 assign n_877 = retime_s6_39_reg_reg_IQ;
 reg retime_s6_40_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_40_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_40_reg_reg_IQ <= sub_561_2_n_22;
     end
 assign n_876 = retime_s6_40_reg_reg_IQ;
 reg retime_s6_41_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_41_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_41_reg_reg_IQ <= sub_561_2_n_86;
     end
 assign n_875 = retime_s6_41_reg_reg_IQ;
 reg retime_s6_42_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_42_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_42_reg_reg_IQ <= n_3621;
     end
 assign n_874 = retime_s6_42_reg_reg_IQ;
 reg retime_s6_43_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_43_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_43_reg_reg_IQ <= sub_561_2_n_27;
     end
 assign n_873 = retime_s6_43_reg_reg_IQ;
 reg retime_s6_44_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_44_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_44_reg_reg_IQ <= n_3371;
     end
 assign n_872 = retime_s6_44_reg_reg_IQ;
 reg retime_s6_45_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_45_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_45_reg_reg_IQ <= n_1941;
     end
 assign n_871 = retime_s6_45_reg_reg_IQ;
 reg retime_s6_46_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_46_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_46_reg_reg_IQ <= n_3372;
     end
 assign n_870 = retime_s6_46_reg_reg_IQ;
 reg retime_s6_47_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_47_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_47_reg_reg_IQ <= n_1943;
     end
 assign n_869 = retime_s6_47_reg_reg_IQ;
 reg retime_s6_48_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_48_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_48_reg_reg_IQ <= n_1942;
     end
 assign n_868 = retime_s6_48_reg_reg_IQ;
 reg retime_s6_49_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_49_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_49_reg_reg_IQ <= n_1944;
     end
 assign n_867 = retime_s6_49_reg_reg_IQ;
 reg retime_s6_50_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_50_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_50_reg_reg_IQ <= n_1921;
     end
 assign n_866 = retime_s6_50_reg_reg_IQ;
 reg retime_s6_51_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_51_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_51_reg_reg_IQ <= n_3374;
     end
 assign n_865 = retime_s6_51_reg_reg_IQ;
 reg retime_s6_52_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_52_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_52_reg_reg_IQ <= n_3376;
     end
 assign n_864 = retime_s6_52_reg_reg_IQ;
 reg retime_s6_53_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_53_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_53_reg_reg_IQ <= sub_561_2_n_14;
     end
 assign n_863 = retime_s6_53_reg_reg_IQ;
 reg retime_s6_54_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_54_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_54_reg_reg_IQ <= sub_561_2_n_42;
     end
 assign n_862 = retime_s6_54_reg_reg_IQ;
 reg retime_s6_55_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_55_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_55_reg_reg_IQ <= n_3378;
     end
 assign n_861 = retime_s6_55_reg_reg_IQ;
 reg retime_s6_56_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_56_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_56_reg_reg_IQ <= n_3379;
     end
 assign n_860 = retime_s6_56_reg_reg_IQ;
 reg retime_s6_57_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_57_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_57_reg_reg_IQ <= sub_561_2_n_9;
     end
 assign n_859 = retime_s6_57_reg_reg_IQ;
 reg retime_s6_58_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_58_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_58_reg_reg_IQ <= sub_561_2_n_20;
     end
 assign n_858 = retime_s6_58_reg_reg_IQ;
 reg retime_s6_59_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_59_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_59_reg_reg_IQ <= sub_561_2_n_39;
     end
 assign n_857 = retime_s6_59_reg_reg_IQ;
 reg retime_s6_60_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_60_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_60_reg_reg_IQ <= n_3381;
     end
 assign n_856 = retime_s6_60_reg_reg_IQ;
 reg retime_s6_61_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_61_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_61_reg_reg_IQ <= n_3377;
     end
 assign n_855 = retime_s6_61_reg_reg_IQ;
 reg retime_s6_62_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_62_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_62_reg_reg_IQ <= n_1945;
     end
 assign n_854 = retime_s6_62_reg_reg_IQ;
 reg retime_s6_65_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_65_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_65_reg_reg_IQ <= n_294;
     end
 assign n_710 = retime_s6_65_reg_reg_IQ;
 reg retime_s6_67_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_67_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_67_reg_reg_IQ <= n_701;
     end
 assign n_700 = retime_s6_67_reg_reg_IQ;
 reg retime_s6_68_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_68_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_68_reg_reg_IQ <= n_689;
     end
 assign n_688 = retime_s6_68_reg_reg_IQ;
 reg retime_s6_69_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_69_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_69_reg_reg_IQ <= n_679;
     end
 assign n_678 = retime_s6_69_reg_reg_IQ;
 reg retime_s6_71_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_71_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_71_reg_reg_IQ <= n_287;
     end
 assign n_672 = retime_s6_71_reg_reg_IQ;
 reg retime_s6_72_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_72_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_72_reg_reg_IQ <= n_666;
     end
 assign n_665 = retime_s6_72_reg_reg_IQ;
 reg retime_s6_73_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_73_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_73_reg_reg_IQ <= n_656;
     end
 assign n_655 = retime_s6_73_reg_reg_IQ;
 reg retime_s6_74_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_74_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_74_reg_reg_IQ <= n_638;
     end
 assign n_637 = retime_s6_74_reg_reg_IQ;
 reg retime_s6_75_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_75_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_75_reg_reg_IQ <= n_624;
     end
 assign n_623 = retime_s6_75_reg_reg_IQ;
 reg retime_s6_76_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_76_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_76_reg_reg_IQ <= n_610;
     end
 assign n_609 = retime_s6_76_reg_reg_IQ;
 reg retime_s6_77_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_77_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_77_reg_reg_IQ <= n_600;
     end
 assign n_599 = retime_s6_77_reg_reg_IQ;
 reg retime_s6_78_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_78_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_78_reg_reg_IQ <= n_590;
     end
 assign n_589 = retime_s6_78_reg_reg_IQ;
 reg retime_s6_79_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_79_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_79_reg_reg_IQ <= n_35;
     end
 assign n_574 = retime_s6_79_reg_reg_IQ;
 reg retime_s6_81_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_81_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_81_reg_reg_IQ <= n_98;
     end
 assign n_572 = retime_s6_81_reg_reg_IQ;
 reg retime_s6_83_reg_reg_IQ;
 wire retime_s6_83_reg_reg_IQN;
 assign retime_s6_83_reg_reg_IQN = !retime_s6_83_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_83_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_83_reg_reg_IQ <= n_284;
     end
 assign n_283 = retime_s6_83_reg_reg_IQN;
 reg retime_s6_84_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_84_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_84_reg_reg_IQ <= n_281;
     end
 assign n_569 = retime_s6_84_reg_reg_IQ;
 reg retime_s6_85_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_85_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_85_reg_reg_IQ <= n_564;
     end
 assign n_563 = retime_s6_85_reg_reg_IQ;
 reg retime_s6_86_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_86_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_86_reg_reg_IQ <= n_554;
     end
 assign n_553 = retime_s6_86_reg_reg_IQ;
 reg retime_s6_87_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_87_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_87_reg_reg_IQ <= n_544;
     end
 assign n_543 = retime_s6_87_reg_reg_IQ;
 reg retime_s6_88_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_88_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_88_reg_reg_IQ <= n_534;
     end
 assign n_533 = retime_s6_88_reg_reg_IQ;
 reg retime_s6_89_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_89_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_89_reg_reg_IQ <= n_523;
     end
 assign n_522 = retime_s6_89_reg_reg_IQ;
 reg retime_s6_93_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_93_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_93_reg_reg_IQ <= n_94;
     end
 assign n_514 = retime_s6_93_reg_reg_IQ;
 reg retime_s6_94_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_94_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_94_reg_reg_IQ <= n_93;
     end
 assign n_513 = retime_s6_94_reg_reg_IQ;
 reg retime_s6_95_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_95_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_95_reg_reg_IQ <= n_278;
     end
 assign n_512 = retime_s6_95_reg_reg_IQ;
 reg retime_s6_100_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_100_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_100_reg_reg_IQ <= n_503;
     end
 assign n_502 = retime_s6_100_reg_reg_IQ;
 reg retime_s6_102_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_102_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_102_reg_reg_IQ <= n_482;
     end
 assign n_481 = retime_s6_102_reg_reg_IQ;
 reg retime_s6_103_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_103_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_103_reg_reg_IQ <= n_472;
     end
 assign n_471 = retime_s6_103_reg_reg_IQ;
 reg retime_s6_104_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_104_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_104_reg_reg_IQ <= n_462;
     end
 assign n_461 = retime_s6_104_reg_reg_IQ;
 reg retime_s6_105_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_105_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_105_reg_reg_IQ <= n_452;
     end
 assign n_451 = retime_s6_105_reg_reg_IQ;
 reg retime_s6_106_reg_reg_IQ;
 wire retime_s6_106_reg_reg_IQN;
 assign retime_s6_106_reg_reg_IQN = !retime_s6_106_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_106_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_106_reg_reg_IQ <= n_273;
     end
 assign n_272 = retime_s6_106_reg_reg_IQN;
 reg retime_s6_107_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_107_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_107_reg_reg_IQ <= n_441;
     end
 assign n_440 = retime_s6_107_reg_reg_IQ;
 reg retime_s6_108_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_108_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_108_reg_reg_IQ <= n_431;
     end
 assign n_430 = retime_s6_108_reg_reg_IQ;
 reg retime_s6_109_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_109_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_109_reg_reg_IQ <= n_421;
     end
 assign n_420 = retime_s6_109_reg_reg_IQ;
 reg retime_s6_110_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_110_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_110_reg_reg_IQ <= n_411;
     end
 assign n_410 = retime_s6_110_reg_reg_IQ;
 reg retime_s6_111_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_111_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_111_reg_reg_IQ <= n_397;
     end
 assign n_396 = retime_s6_111_reg_reg_IQ;
 reg retime_s6_112_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_112_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_112_reg_reg_IQ <= n_387;
     end
 assign n_386 = retime_s6_112_reg_reg_IQ;
 reg retime_s6_117_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_117_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_117_reg_reg_IQ <= n_372;
     end
 assign n_371 = retime_s6_117_reg_reg_IQ;
 reg retime_s6_119_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_119_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_119_reg_reg_IQ <= n_361;
     end
 assign n_360 = retime_s6_119_reg_reg_IQ;
 reg retime_s6_120_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_120_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_120_reg_reg_IQ <= n_351;
     end
 assign n_350 = retime_s6_120_reg_reg_IQ;
 reg retime_s6_122_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_122_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_122_reg_reg_IQ <= n_340;
     end
 assign n_339 = retime_s6_122_reg_reg_IQ;
 reg retime_s7_3_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_3_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_3_reg_reg_IQ <= n_1110;
     end
 assign n_1109 = retime_s7_3_reg_reg_IQ;
 reg retime_s7_4_reg_reg_IQ;
 wire retime_s7_4_reg_reg_IQN;
 assign retime_s7_4_reg_reg_IQN = !retime_s7_4_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_4_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_4_reg_reg_IQ <= n_300;
     end
 assign n_938 = retime_s7_4_reg_reg_IQN;
 reg retime_s7_5_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_5_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_5_reg_reg_IQ <= n_3448;
     end
 assign n_937 = retime_s7_5_reg_reg_IQ;
 reg retime_s7_6_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_6_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_6_reg_reg_IQ <= n_3430;
     end
 assign n_936 = retime_s7_6_reg_reg_IQ;
 reg retime_s7_7_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_7_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_7_reg_reg_IQ <= n_3441;
     end
 assign n_935 = retime_s7_7_reg_reg_IQ;
 reg retime_s7_8_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_8_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_8_reg_reg_IQ <= n_3443;
     end
 assign n_934 = retime_s7_8_reg_reg_IQ;
 reg retime_s7_9_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_9_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_9_reg_reg_IQ <= n_3432;
     end
 assign n_933 = retime_s7_9_reg_reg_IQ;
 reg retime_s7_10_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_10_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_10_reg_reg_IQ <= n_3433;
     end
 assign n_932 = retime_s7_10_reg_reg_IQ;
 reg retime_s7_11_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_11_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_11_reg_reg_IQ <= n_3436;
     end
 assign n_931 = retime_s7_11_reg_reg_IQ;
 reg retime_s7_12_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_12_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_12_reg_reg_IQ <= n_3440;
     end
 assign n_930 = retime_s7_12_reg_reg_IQ;
 reg retime_s7_13_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_13_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_13_reg_reg_IQ <= n_3438;
     end
 assign n_929 = retime_s7_13_reg_reg_IQ;
 reg retime_s7_14_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_14_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_14_reg_reg_IQ <= n_3442;
     end
 assign n_928 = retime_s7_14_reg_reg_IQ;
 reg retime_s7_15_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_15_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_15_reg_reg_IQ <= n_3444;
     end
 assign n_927 = retime_s7_15_reg_reg_IQ;
 reg retime_s7_16_reg_reg_IQ;
 wire retime_s7_16_reg_reg_IQN;
 assign retime_s7_16_reg_reg_IQN = !retime_s7_16_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_16_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_16_reg_reg_IQ <= n_3693;
     end
 assign n_926 = retime_s7_16_reg_reg_IQN;
 reg retime_s7_17_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_17_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_17_reg_reg_IQ <= n_3431;
     end
 assign n_925 = retime_s7_17_reg_reg_IQ;
 reg retime_s7_18_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_18_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_18_reg_reg_IQ <= n_3429;
     end
 assign n_924 = retime_s7_18_reg_reg_IQ;
 reg retime_s7_19_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_19_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_19_reg_reg_IQ <= n_3428;
     end
 assign n_923 = retime_s7_19_reg_reg_IQ;
 reg retime_s7_20_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_20_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_20_reg_reg_IQ <= n_3434;
     end
 assign n_922 = retime_s7_20_reg_reg_IQ;
 reg retime_s7_21_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_21_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_21_reg_reg_IQ <= n_2897;
     end
 assign n_921 = retime_s7_21_reg_reg_IQ;
 reg retime_s7_22_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_22_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_22_reg_reg_IQ <= n_3446;
     end
 assign n_920 = retime_s7_22_reg_reg_IQ;
 reg retime_s7_23_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_23_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_23_reg_reg_IQ <= n_3437;
     end
 assign n_919 = retime_s7_23_reg_reg_IQ;
 reg retime_s7_24_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_24_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_24_reg_reg_IQ <= n_3445;
     end
 assign n_918 = retime_s7_24_reg_reg_IQ;
 reg retime_s7_25_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_25_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_25_reg_reg_IQ <= n_3447;
     end
 assign n_917 = retime_s7_25_reg_reg_IQ;
 reg retime_s7_26_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_26_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_26_reg_reg_IQ <= n_3427;
     end
 assign n_916 = retime_s7_26_reg_reg_IQ;
 reg retime_s7_27_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_27_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_27_reg_reg_IQ <= n_3435;
     end
 assign n_915 = retime_s7_27_reg_reg_IQ;
 reg retime_s7_28_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_28_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_28_reg_reg_IQ <= n_3439;
     end
 assign n_914 = retime_s7_28_reg_reg_IQ;
 reg retime_s7_29_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_29_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_29_reg_reg_IQ <= n_3409;
     end
 assign n_913 = retime_s7_29_reg_reg_IQ;
 reg retime_s7_30_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_30_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_30_reg_reg_IQ <= n_145;
     end
 assign n_720 = retime_s7_30_reg_reg_IQ;
 reg retime_s7_31_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_31_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_31_reg_reg_IQ <= n_142;
     end
 assign n_719 = retime_s7_31_reg_reg_IQ;
 reg retime_s7_32_reg_reg_IQ;
 wire retime_s7_32_reg_reg_IQN;
 assign retime_s7_32_reg_reg_IQN = !retime_s7_32_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_32_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_32_reg_reg_IQ <= n_146;
     end
 assign n_291 = retime_s7_32_reg_reg_IQN;
 reg retime_s7_33_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_33_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_33_reg_reg_IQ <= n_700;
     end
 assign n_699 = retime_s7_33_reg_reg_IQ;
 reg retime_s7_34_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_34_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_34_reg_reg_IQ <= n_688;
     end
 assign n_687 = retime_s7_34_reg_reg_IQ;
 reg retime_s7_35_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_35_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_35_reg_reg_IQ <= n_678;
     end
 assign n_677 = retime_s7_35_reg_reg_IQ;
 reg retime_s7_37_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_37_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_37_reg_reg_IQ <= n_665;
     end
 assign n_664 = retime_s7_37_reg_reg_IQ;
 reg retime_s7_38_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_38_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_38_reg_reg_IQ <= n_655;
     end
 assign n_654 = retime_s7_38_reg_reg_IQ;
 reg retime_s7_39_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_39_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_39_reg_reg_IQ <= n_637;
     end
 assign n_636 = retime_s7_39_reg_reg_IQ;
 reg retime_s7_40_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_40_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_40_reg_reg_IQ <= n_623;
     end
 assign n_622 = retime_s7_40_reg_reg_IQ;
 reg retime_s7_41_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_41_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_41_reg_reg_IQ <= n_609;
     end
 assign n_608 = retime_s7_41_reg_reg_IQ;
 reg retime_s7_42_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_42_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_42_reg_reg_IQ <= n_599;
     end
 assign n_598 = retime_s7_42_reg_reg_IQ;
 reg retime_s7_43_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_43_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_43_reg_reg_IQ <= n_589;
     end
 assign n_588 = retime_s7_43_reg_reg_IQ;
 reg retime_s7_45_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_45_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_45_reg_reg_IQ <= n_74;
     end
 assign n_571 = retime_s7_45_reg_reg_IQ;
 reg retime_s7_46_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_46_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_46_reg_reg_IQ <= n_283;
     end
 assign n_282 = retime_s7_46_reg_reg_IQ;
 reg retime_s7_47_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_47_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_47_reg_reg_IQ <= n_563;
     end
 assign n_562 = retime_s7_47_reg_reg_IQ;
 reg retime_s7_48_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_48_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_48_reg_reg_IQ <= n_553;
     end
 assign n_552 = retime_s7_48_reg_reg_IQ;
 reg retime_s7_49_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_49_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_49_reg_reg_IQ <= n_543;
     end
 assign n_542 = retime_s7_49_reg_reg_IQ;
 reg retime_s7_50_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_50_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_50_reg_reg_IQ <= n_533;
     end
 assign n_532 = retime_s7_50_reg_reg_IQ;
 reg retime_s7_51_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_51_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_51_reg_reg_IQ <= n_522;
     end
 assign n_521 = retime_s7_51_reg_reg_IQ;
 reg retime_s7_54_reg_reg_IQ;
 wire retime_s7_54_reg_reg_IQN;
 assign retime_s7_54_reg_reg_IQN = !retime_s7_54_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_54_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_54_reg_reg_IQ <= n_163;
     end
 assign n_279 = retime_s7_54_reg_reg_IQN;
 reg retime_s7_58_reg_reg_IQ;
 wire retime_s7_58_reg_reg_IQN;
 assign retime_s7_58_reg_reg_IQN = !retime_s7_58_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_58_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_58_reg_reg_IQ <= n_21;
     end
 assign n_276 = retime_s7_58_reg_reg_IQN;
 reg retime_s7_59_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_59_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_59_reg_reg_IQ <= n_502;
     end
 assign n_501 = retime_s7_59_reg_reg_IQ;
 reg retime_s7_61_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_61_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_61_reg_reg_IQ <= n_481;
     end
 assign n_480 = retime_s7_61_reg_reg_IQ;
 reg retime_s7_62_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_62_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_62_reg_reg_IQ <= n_471;
     end
 assign n_470 = retime_s7_62_reg_reg_IQ;
 reg retime_s7_63_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_63_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_63_reg_reg_IQ <= n_461;
     end
 assign n_460 = retime_s7_63_reg_reg_IQ;
 reg retime_s7_64_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_64_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_64_reg_reg_IQ <= n_451;
     end
 assign n_450 = retime_s7_64_reg_reg_IQ;
 reg retime_s7_65_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_65_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_65_reg_reg_IQ <= n_272;
     end
 assign n_446 = retime_s7_65_reg_reg_IQ;
 reg retime_s7_66_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_66_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_66_reg_reg_IQ <= n_440;
     end
 assign n_439 = retime_s7_66_reg_reg_IQ;
 reg retime_s7_67_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_67_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_67_reg_reg_IQ <= n_430;
     end
 assign n_429 = retime_s7_67_reg_reg_IQ;
 reg retime_s7_68_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_68_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_68_reg_reg_IQ <= n_420;
     end
 assign n_419 = retime_s7_68_reg_reg_IQ;
 reg retime_s7_69_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_69_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_69_reg_reg_IQ <= n_410;
     end
 assign n_409 = retime_s7_69_reg_reg_IQ;
 reg retime_s7_70_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_70_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_70_reg_reg_IQ <= n_396;
     end
 assign n_395 = retime_s7_70_reg_reg_IQ;
 reg retime_s7_71_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_71_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_71_reg_reg_IQ <= n_386;
     end
 assign n_385 = retime_s7_71_reg_reg_IQ;
 reg retime_s7_73_reg_reg_IQ;
 wire retime_s7_73_reg_reg_IQN;
 assign retime_s7_73_reg_reg_IQN = !retime_s7_73_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_73_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_73_reg_reg_IQ <= n_70;
     end
 assign n_270 = retime_s7_73_reg_reg_IQN;
 reg retime_s7_74_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_74_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_74_reg_reg_IQ <= n_177;
     end
 assign n_378 = retime_s7_74_reg_reg_IQ;
 reg retime_s7_75_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_75_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_75_reg_reg_IQ <= n_180;
     end
 assign n_377 = retime_s7_75_reg_reg_IQ;
 reg retime_s7_76_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_76_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_76_reg_reg_IQ <= n_371;
     end
 assign n_370 = retime_s7_76_reg_reg_IQ;
 reg retime_s7_78_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_78_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_78_reg_reg_IQ <= n_360;
     end
 assign n_359 = retime_s7_78_reg_reg_IQ;
 reg retime_s7_79_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_79_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_79_reg_reg_IQ <= n_350;
     end
 assign n_349 = retime_s7_79_reg_reg_IQ;
 reg retime_s7_80_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_80_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_80_reg_reg_IQ <= n_104;
     end
 assign n_345 = retime_s7_80_reg_reg_IQ;
 reg retime_s7_81_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_81_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_81_reg_reg_IQ <= n_339;
     end
 assign n_338 = retime_s7_81_reg_reg_IQ;
 reg retime_s8_3_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_3_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_3_reg_reg_IQ <= n_1109;
     end
 assign n_1108 = retime_s8_3_reg_reg_IQ;
 reg retime_s8_4_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_4_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_4_reg_reg_IQ <= sub_656_2_n_52;
     end
 assign n_1015 = retime_s8_4_reg_reg_IQ;
 reg retime_s8_5_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_5_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_5_reg_reg_IQ <= n_3487;
     end
 assign n_1014 = retime_s8_5_reg_reg_IQ;
 reg retime_s8_6_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_6_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_6_reg_reg_IQ <= sub_656_2_n_68;
     end
 assign n_1013 = retime_s8_6_reg_reg_IQ;
 reg retime_s8_7_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_7_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_7_reg_reg_IQ <= n_3480;
     end
 assign n_1012 = retime_s8_7_reg_reg_IQ;
 reg retime_s8_8_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_8_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_8_reg_reg_IQ <= sub_656_2_n_83;
     end
 assign n_1011 = retime_s8_8_reg_reg_IQ;
 reg retime_s8_9_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_9_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_9_reg_reg_IQ <= sub_656_2_n_118;
     end
 assign n_1010 = retime_s8_9_reg_reg_IQ;
 reg retime_s8_10_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_10_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_10_reg_reg_IQ <= n_3478;
     end
 assign n_1009 = retime_s8_10_reg_reg_IQ;
 reg retime_s8_11_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_11_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_11_reg_reg_IQ <= n_3475;
     end
 assign n_1008 = retime_s8_11_reg_reg_IQ;
 reg retime_s8_12_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_12_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_12_reg_reg_IQ <= n_3484;
     end
 assign n_1007 = retime_s8_12_reg_reg_IQ;
 reg retime_s8_13_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_13_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_13_reg_reg_IQ <= n_3473;
     end
 assign n_1006 = retime_s8_13_reg_reg_IQ;
 reg retime_s8_14_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_14_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_14_reg_reg_IQ <= sub_656_2_n_65;
     end
 assign n_1005 = retime_s8_14_reg_reg_IQ;
 reg retime_s8_15_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_15_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_15_reg_reg_IQ <= sub_656_2_n_136;
     end
 assign n_1004 = retime_s8_15_reg_reg_IQ;
 reg retime_s8_16_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_16_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_16_reg_reg_IQ <= n_2189;
     end
 assign n_1003 = retime_s8_16_reg_reg_IQ;
 reg retime_s8_17_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_17_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_17_reg_reg_IQ <= n_3711;
     end
 assign n_1002 = retime_s8_17_reg_reg_IQ;
 reg retime_s8_18_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_18_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_18_reg_reg_IQ <= n_2187;
     end
 assign n_1001 = retime_s8_18_reg_reg_IQ;
 reg retime_s8_19_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_19_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_19_reg_reg_IQ <= n_2188;
     end
 assign n_1000 = retime_s8_19_reg_reg_IQ;
 reg retime_s8_20_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_20_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_20_reg_reg_IQ <= sub_656_2_n_126;
     end
 assign n_999 = retime_s8_20_reg_reg_IQ;
 reg retime_s8_21_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_21_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_21_reg_reg_IQ <= sub_656_2_n_70;
     end
 assign n_998 = retime_s8_21_reg_reg_IQ;
 reg retime_s8_22_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_22_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_22_reg_reg_IQ <= sub_656_2_n_111;
     end
 assign n_997 = retime_s8_22_reg_reg_IQ;
 reg retime_s8_23_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_23_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_23_reg_reg_IQ <= sub_656_2_n_164;
     end
 assign n_996 = retime_s8_23_reg_reg_IQ;
 reg retime_s8_24_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_24_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_24_reg_reg_IQ <= sub_656_2_n_168;
     end
 assign n_995 = retime_s8_24_reg_reg_IQ;
 reg retime_s8_25_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_25_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_25_reg_reg_IQ <= n_3476;
     end
 assign n_994 = retime_s8_25_reg_reg_IQ;
 reg retime_s8_26_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_26_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_26_reg_reg_IQ <= sub_656_2_n_88;
     end
 assign n_993 = retime_s8_26_reg_reg_IQ;
 reg retime_s8_27_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_27_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_27_reg_reg_IQ <= n_3470;
     end
 assign n_992 = retime_s8_27_reg_reg_IQ;
 reg retime_s8_28_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_28_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_28_reg_reg_IQ <= sub_656_2_n_19;
     end
 assign n_991 = retime_s8_28_reg_reg_IQ;
 reg retime_s8_29_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_29_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_29_reg_reg_IQ <= sub_656_2_n_134;
     end
 assign n_990 = retime_s8_29_reg_reg_IQ;
 reg retime_s8_30_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_30_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_30_reg_reg_IQ <= sub_656_2_n_147;
     end
 assign n_989 = retime_s8_30_reg_reg_IQ;
 reg retime_s8_31_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_31_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_31_reg_reg_IQ <= n_3489;
     end
 assign n_988 = retime_s8_31_reg_reg_IQ;
 reg retime_s8_32_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_32_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_32_reg_reg_IQ <= sub_656_2_n_108;
     end
 assign n_987 = retime_s8_32_reg_reg_IQ;
 reg retime_s8_33_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_33_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_33_reg_reg_IQ <= sub_656_2_n_127;
     end
 assign n_986 = retime_s8_33_reg_reg_IQ;
 reg retime_s8_34_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_34_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_34_reg_reg_IQ <= n_3481;
     end
 assign n_985 = retime_s8_34_reg_reg_IQ;
 reg retime_s8_35_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_35_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_35_reg_reg_IQ <= n_3479;
     end
 assign n_984 = retime_s8_35_reg_reg_IQ;
 reg retime_s8_36_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_36_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_36_reg_reg_IQ <= sub_656_2_n_72;
     end
 assign n_983 = retime_s8_36_reg_reg_IQ;
 reg retime_s8_37_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_37_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_37_reg_reg_IQ <= sub_656_2_n_75;
     end
 assign n_982 = retime_s8_37_reg_reg_IQ;
 reg retime_s8_38_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_38_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_38_reg_reg_IQ <= n_3474;
     end
 assign n_981 = retime_s8_38_reg_reg_IQ;
 reg retime_s8_39_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_39_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_39_reg_reg_IQ <= sub_656_2_n_9;
     end
 assign n_980 = retime_s8_39_reg_reg_IQ;
 reg retime_s8_40_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_40_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_40_reg_reg_IQ <= sub_656_2_n_105;
     end
 assign n_979 = retime_s8_40_reg_reg_IQ;
 reg retime_s8_41_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_41_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_41_reg_reg_IQ <= sub_656_2_n_132;
     end
 assign n_978 = retime_s8_41_reg_reg_IQ;
 reg retime_s8_42_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_42_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_42_reg_reg_IQ <= n_3677;
     end
 assign n_977 = retime_s8_42_reg_reg_IQ;
 reg retime_s8_43_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_43_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_43_reg_reg_IQ <= sub_656_2_n_29;
     end
 assign n_976 = retime_s8_43_reg_reg_IQ;
 reg retime_s8_44_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_44_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_44_reg_reg_IQ <= n_3482;
     end
 assign n_975 = retime_s8_44_reg_reg_IQ;
 reg retime_s8_45_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_45_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_45_reg_reg_IQ <= sub_656_2_n_94;
     end
 assign n_974 = retime_s8_45_reg_reg_IQ;
 reg retime_s8_46_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_46_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_46_reg_reg_IQ <= sub_656_2_n_120;
     end
 assign n_973 = retime_s8_46_reg_reg_IQ;
 reg retime_s8_47_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_47_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_47_reg_reg_IQ <= n_3488;
     end
 assign n_972 = retime_s8_47_reg_reg_IQ;
 reg retime_s8_48_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_48_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_48_reg_reg_IQ <= n_3471;
     end
 assign n_971 = retime_s8_48_reg_reg_IQ;
 reg retime_s8_49_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_49_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_49_reg_reg_IQ <= sub_656_2_n_91;
     end
 assign n_970 = retime_s8_49_reg_reg_IQ;
 reg retime_s8_50_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_50_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_50_reg_reg_IQ <= n_2190;
     end
 assign n_969 = retime_s8_50_reg_reg_IQ;
 reg retime_s8_51_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_51_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_51_reg_reg_IQ <= n_2191;
     end
 assign n_968 = retime_s8_51_reg_reg_IQ;
 reg retime_s8_52_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_52_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_52_reg_reg_IQ <= sub_656_2_n_143;
     end
 assign n_967 = retime_s8_52_reg_reg_IQ;
 reg retime_s8_53_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_53_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_53_reg_reg_IQ <= sub_656_2_n_66;
     end
 assign n_966 = retime_s8_53_reg_reg_IQ;
 reg retime_s8_54_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_54_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_54_reg_reg_IQ <= sub_656_2_n_124;
     end
 assign n_965 = retime_s8_54_reg_reg_IQ;
 reg retime_s8_55_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_55_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_55_reg_reg_IQ <= n_3472;
     end
 assign n_964 = retime_s8_55_reg_reg_IQ;
 reg retime_s8_56_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_56_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_56_reg_reg_IQ <= n_3483;
     end
 assign n_963 = retime_s8_56_reg_reg_IQ;
 reg retime_s8_57_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_57_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_57_reg_reg_IQ <= sub_656_2_n_11;
     end
 assign n_962 = retime_s8_57_reg_reg_IQ;
 reg retime_s8_58_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_58_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_58_reg_reg_IQ <= n_3063;
     end
 assign n_961 = retime_s8_58_reg_reg_IQ;
 reg retime_s8_59_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_59_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_59_reg_reg_IQ <= n_2195;
     end
 assign n_960 = retime_s8_59_reg_reg_IQ;
 reg retime_s8_60_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_60_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_60_reg_reg_IQ <= sub_656_2_n_55;
     end
 assign n_959 = retime_s8_60_reg_reg_IQ;
 reg retime_s8_61_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_61_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_61_reg_reg_IQ <= n_2194;
     end
 assign n_958 = retime_s8_61_reg_reg_IQ;
 reg retime_s8_62_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_62_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_62_reg_reg_IQ <= n_2193;
     end
 assign n_957 = retime_s8_62_reg_reg_IQ;
 reg retime_s8_63_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_63_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_63_reg_reg_IQ <= n_2192;
     end
 assign n_956 = retime_s8_63_reg_reg_IQ;
 reg retime_s8_64_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_64_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_64_reg_reg_IQ <= n_2160;
     end
 assign n_955 = retime_s8_64_reg_reg_IQ;
 reg retime_s8_65_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_65_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_65_reg_reg_IQ <= n_3486;
     end
 assign n_954 = retime_s8_65_reg_reg_IQ;
 reg retime_s8_66_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_66_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_66_reg_reg_IQ <= sub_656_2_n_89;
     end
 assign n_953 = retime_s8_66_reg_reg_IQ;
 reg retime_s8_67_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_67_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_67_reg_reg_IQ <= sub_656_2_n_123;
     end
 assign n_952 = retime_s8_67_reg_reg_IQ;
 reg retime_s8_68_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_68_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_68_reg_reg_IQ <= sub_656_2_n_100;
     end
 assign n_951 = retime_s8_68_reg_reg_IQ;
 reg retime_s8_69_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_69_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_69_reg_reg_IQ <= n_2166;
     end
 assign n_950 = retime_s8_69_reg_reg_IQ;
 reg retime_s8_70_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_70_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_70_reg_reg_IQ <= n_3491;
     end
 assign n_949 = retime_s8_70_reg_reg_IQ;
 reg retime_s8_71_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_71_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_71_reg_reg_IQ <= n_3062;
     end
 assign n_948 = retime_s8_71_reg_reg_IQ;
 reg retime_s8_72_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_72_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_72_reg_reg_IQ <= sub_656_2_n_49;
     end
 assign n_947 = retime_s8_72_reg_reg_IQ;
 reg retime_s8_73_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_73_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_73_reg_reg_IQ <= sub_656_2_n_47;
     end
 assign n_946 = retime_s8_73_reg_reg_IQ;
 reg retime_s8_74_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_74_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_74_reg_reg_IQ <= n_3477;
     end
 assign n_945 = retime_s8_74_reg_reg_IQ;
 reg retime_s8_75_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_75_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_75_reg_reg_IQ <= sub_656_2_n_56;
     end
 assign n_944 = retime_s8_75_reg_reg_IQ;
 reg retime_s8_76_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_76_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_76_reg_reg_IQ <= sub_656_2_n_71;
     end
 assign n_943 = retime_s8_76_reg_reg_IQ;
 reg retime_s8_77_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_77_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_77_reg_reg_IQ <= sub_656_2_n_54;
     end
 assign n_942 = retime_s8_77_reg_reg_IQ;
 reg retime_s8_78_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_78_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_78_reg_reg_IQ <= n_3490;
     end
 assign n_941 = retime_s8_78_reg_reg_IQ;
 reg retime_s8_79_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_79_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_79_reg_reg_IQ <= sub_656_2_n_43;
     end
 assign n_940 = retime_s8_79_reg_reg_IQ;
 reg retime_s8_80_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_80_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_80_reg_reg_IQ <= n_3485;
     end
 assign n_939 = retime_s8_80_reg_reg_IQ;
 reg retime_s8_81_reg_reg_IQ;
 wire retime_s8_81_reg_reg_IQN;
 assign retime_s8_81_reg_reg_IQN = !retime_s8_81_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_81_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_81_reg_reg_IQ <= n_291;
     end
 assign n_290 = retime_s8_81_reg_reg_IQN;
 reg retime_s8_82_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_82_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_82_reg_reg_IQ <= n_699;
     end
 assign n_698 = retime_s8_82_reg_reg_IQ;
 reg retime_s8_83_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_83_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_83_reg_reg_IQ <= n_687;
     end
 assign n_686 = retime_s8_83_reg_reg_IQ;
 reg retime_s8_84_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_84_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_84_reg_reg_IQ <= n_677;
     end
 assign n_676 = retime_s8_84_reg_reg_IQ;
 reg retime_s8_86_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_86_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_86_reg_reg_IQ <= n_664;
     end
 assign n_663 = retime_s8_86_reg_reg_IQ;
 reg retime_s8_87_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_87_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_87_reg_reg_IQ <= n_654;
     end
 assign n_653 = retime_s8_87_reg_reg_IQ;
 reg retime_s8_88_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_88_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_88_reg_reg_IQ <= n_636;
     end
 assign n_635 = retime_s8_88_reg_reg_IQ;
 reg retime_s8_89_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_89_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_89_reg_reg_IQ <= n_622;
     end
 assign n_621 = retime_s8_89_reg_reg_IQ;
 reg retime_s8_90_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_90_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_90_reg_reg_IQ <= n_608;
     end
 assign n_607 = retime_s8_90_reg_reg_IQ;
 reg retime_s8_91_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_91_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_91_reg_reg_IQ <= n_598;
     end
 assign n_597 = retime_s8_91_reg_reg_IQ;
 reg retime_s8_92_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_92_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_92_reg_reg_IQ <= n_588;
     end
 assign n_587 = retime_s8_92_reg_reg_IQ;
 reg retime_s8_93_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_93_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_93_reg_reg_IQ <= n_58;
     end
 assign n_573 = retime_s8_93_reg_reg_IQ;
 reg retime_s8_94_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_94_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_94_reg_reg_IQ <= n_282;
     end
 assign n_570 = retime_s8_94_reg_reg_IQ;
 reg retime_s8_95_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_95_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_95_reg_reg_IQ <= n_562;
     end
 assign n_561 = retime_s8_95_reg_reg_IQ;
 reg retime_s8_96_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_96_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_96_reg_reg_IQ <= n_552;
     end
 assign n_551 = retime_s8_96_reg_reg_IQ;
 reg retime_s8_97_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_97_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_97_reg_reg_IQ <= n_542;
     end
 assign n_541 = retime_s8_97_reg_reg_IQ;
 reg retime_s8_98_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_98_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_98_reg_reg_IQ <= n_532;
     end
 assign n_531 = retime_s8_98_reg_reg_IQ;
 reg retime_s8_99_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_99_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_99_reg_reg_IQ <= n_521;
     end
 assign n_520 = retime_s8_99_reg_reg_IQ;
 reg retime_s8_100_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_100_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_100_reg_reg_IQ <= n_133;
     end
 assign n_517 = retime_s8_100_reg_reg_IQ;
 reg retime_s8_101_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_101_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_101_reg_reg_IQ <= n_57;
     end
 assign n_516 = retime_s8_101_reg_reg_IQ;
 reg retime_s8_102_reg_reg_IQ;
 wire retime_s8_102_reg_reg_IQN;
 assign retime_s8_102_reg_reg_IQN = !retime_s8_102_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_102_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_102_reg_reg_IQ <= n_279;
     end
 assign n_515 = retime_s8_102_reg_reg_IQN;
 reg retime_s8_106_reg_reg_IQ;
 wire retime_s8_106_reg_reg_IQN;
 assign retime_s8_106_reg_reg_IQN = !retime_s8_106_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_106_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_106_reg_reg_IQ <= n_276;
     end
 assign n_275 = retime_s8_106_reg_reg_IQN;
 reg retime_s8_107_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_107_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_107_reg_reg_IQ <= n_501;
     end
 assign n_500 = retime_s8_107_reg_reg_IQ;
 reg retime_s8_109_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_109_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_109_reg_reg_IQ <= n_480;
     end
 assign n_479 = retime_s8_109_reg_reg_IQ;
 reg retime_s8_110_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_110_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_110_reg_reg_IQ <= n_470;
     end
 assign n_469 = retime_s8_110_reg_reg_IQ;
 reg retime_s8_111_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_111_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_111_reg_reg_IQ <= n_460;
     end
 assign n_459 = retime_s8_111_reg_reg_IQ;
 reg retime_s8_112_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_112_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_112_reg_reg_IQ <= n_450;
     end
 assign n_449 = retime_s8_112_reg_reg_IQ;
 reg retime_s8_113_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_113_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_113_reg_reg_IQ <= n_439;
     end
 assign n_438 = retime_s8_113_reg_reg_IQ;
 reg retime_s8_114_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_114_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_114_reg_reg_IQ <= n_429;
     end
 assign n_428 = retime_s8_114_reg_reg_IQ;
 reg retime_s8_115_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_115_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_115_reg_reg_IQ <= n_419;
     end
 assign n_418 = retime_s8_115_reg_reg_IQ;
 reg retime_s8_116_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_116_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_116_reg_reg_IQ <= n_409;
     end
 assign n_408 = retime_s8_116_reg_reg_IQ;
 reg retime_s8_117_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_117_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_117_reg_reg_IQ <= n_395;
     end
 assign n_394 = retime_s8_117_reg_reg_IQ;
 reg retime_s8_118_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_118_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_118_reg_reg_IQ <= n_385;
     end
 assign n_384 = retime_s8_118_reg_reg_IQ;
 reg retime_s8_119_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_119_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_119_reg_reg_IQ <= n_51;
     end
 assign n_380 = retime_s8_119_reg_reg_IQ;
 reg retime_s8_120_reg_reg_IQ;
 wire retime_s8_120_reg_reg_IQN;
 assign retime_s8_120_reg_reg_IQN = !retime_s8_120_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_120_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_120_reg_reg_IQ <= n_270;
     end
 assign n_379 = retime_s8_120_reg_reg_IQN;
 reg retime_s8_121_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_121_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_121_reg_reg_IQ <= n_370;
     end
 assign n_369 = retime_s8_121_reg_reg_IQ;
 reg retime_s8_122_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_122_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_122_reg_reg_IQ <= n_49;
     end
 assign n_366 = retime_s8_122_reg_reg_IQ;
 reg retime_s8_123_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_123_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_123_reg_reg_IQ <= n_359;
     end
 assign n_358 = retime_s8_123_reg_reg_IQ;
 reg retime_s8_124_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_124_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_124_reg_reg_IQ <= n_349;
     end
 assign n_348 = retime_s8_124_reg_reg_IQ;
 reg retime_s8_125_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_125_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_125_reg_reg_IQ <= n_338;
     end
 assign n_337 = retime_s8_125_reg_reg_IQ;
 reg retime_s9_3_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_3_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_3_reg_reg_IQ <= n_1108;
     end
 assign n_1107 = retime_s9_3_reg_reg_IQ;
 reg retime_s9_4_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_4_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_4_reg_reg_IQ <= n_2254;
     end
 assign n_1047 = retime_s9_4_reg_reg_IQ;
 reg retime_s9_5_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_5_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_5_reg_reg_IQ <= n_2283;
     end
 assign n_1046 = retime_s9_5_reg_reg_IQ;
 reg retime_s9_6_reg_reg_IQ;
 wire retime_s9_6_reg_reg_IQN;
 assign retime_s9_6_reg_reg_IQN = !retime_s9_6_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_6_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_6_reg_reg_IQ <= n_301;
     end
 assign n_1045 = retime_s9_6_reg_reg_IQN;
 reg retime_s9_7_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_7_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_7_reg_reg_IQ <= n_2336;
     end
 assign n_1044 = retime_s9_7_reg_reg_IQ;
 reg retime_s9_8_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_8_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_8_reg_reg_IQ <= n_2323;
     end
 assign n_1043 = retime_s9_8_reg_reg_IQ;
 reg retime_s9_9_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_9_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_9_reg_reg_IQ <= n_2335;
     end
 assign n_1042 = retime_s9_9_reg_reg_IQ;
 reg retime_s9_10_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_10_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_10_reg_reg_IQ <= n_2334;
     end
 assign n_1041 = retime_s9_10_reg_reg_IQ;
 reg retime_s9_11_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_11_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_11_reg_reg_IQ <= n_2332;
     end
 assign n_1040 = retime_s9_11_reg_reg_IQ;
 reg retime_s9_12_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_12_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_12_reg_reg_IQ <= n_2333;
     end
 assign n_1039 = retime_s9_12_reg_reg_IQ;
 reg retime_s9_13_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_13_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_13_reg_reg_IQ <= n_2322;
     end
 assign n_1038 = retime_s9_13_reg_reg_IQ;
 reg retime_s9_14_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_14_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_14_reg_reg_IQ <= n_2320;
     end
 assign n_1037 = retime_s9_14_reg_reg_IQ;
 reg retime_s9_15_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_15_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_15_reg_reg_IQ <= n_2329;
     end
 assign n_1036 = retime_s9_15_reg_reg_IQ;
 reg retime_s9_16_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_16_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_16_reg_reg_IQ <= n_2319;
     end
 assign n_1035 = retime_s9_16_reg_reg_IQ;
 reg retime_s9_17_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_17_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_17_reg_reg_IQ <= n_2330;
     end
 assign n_1034 = retime_s9_17_reg_reg_IQ;
 reg retime_s9_18_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_18_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_18_reg_reg_IQ <= n_2331;
     end
 assign n_1033 = retime_s9_18_reg_reg_IQ;
 reg retime_s9_19_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_19_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_19_reg_reg_IQ <= n_2311;
     end
 assign n_1032 = retime_s9_19_reg_reg_IQ;
 reg retime_s9_20_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_20_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_20_reg_reg_IQ <= n_2327;
     end
 assign n_1031 = retime_s9_20_reg_reg_IQ;
 reg retime_s9_21_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_21_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_21_reg_reg_IQ <= n_2315;
     end
 assign n_1030 = retime_s9_21_reg_reg_IQ;
 reg retime_s9_22_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_22_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_22_reg_reg_IQ <= n_2326;
     end
 assign n_1029 = retime_s9_22_reg_reg_IQ;
 reg retime_s9_23_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_23_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_23_reg_reg_IQ <= n_2325;
     end
 assign n_1028 = retime_s9_23_reg_reg_IQ;
 reg retime_s9_24_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_24_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_24_reg_reg_IQ <= n_2321;
     end
 assign n_1027 = retime_s9_24_reg_reg_IQ;
 reg retime_s9_25_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_25_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_25_reg_reg_IQ <= n_2339;
     end
 assign n_1026 = retime_s9_25_reg_reg_IQ;
 reg retime_s9_26_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_26_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_26_reg_reg_IQ <= n_2338;
     end
 assign n_1025 = retime_s9_26_reg_reg_IQ;
 reg retime_s9_27_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_27_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_27_reg_reg_IQ <= n_301;
     end
 assign n_1024 = retime_s9_27_reg_reg_IQ;
 reg retime_s9_28_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_28_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_28_reg_reg_IQ <= n_2328;
     end
 assign n_1023 = retime_s9_28_reg_reg_IQ;
 reg retime_s9_29_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_29_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_29_reg_reg_IQ <= n_2314;
     end
 assign n_1022 = retime_s9_29_reg_reg_IQ;
 reg retime_s9_30_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_30_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_30_reg_reg_IQ <= n_2337;
     end
 assign n_1021 = retime_s9_30_reg_reg_IQ;
 reg retime_s9_31_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_31_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_31_reg_reg_IQ <= n_2317;
     end
 assign n_1020 = retime_s9_31_reg_reg_IQ;
 reg retime_s9_32_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_32_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_32_reg_reg_IQ <= n_2318;
     end
 assign n_1019 = retime_s9_32_reg_reg_IQ;
 reg retime_s9_33_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_33_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_33_reg_reg_IQ <= n_2313;
     end
 assign n_1018 = retime_s9_33_reg_reg_IQ;
 reg retime_s9_34_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_34_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_34_reg_reg_IQ <= n_2324;
     end
 assign n_1017 = retime_s9_34_reg_reg_IQ;
 reg retime_s9_35_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_35_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_35_reg_reg_IQ <= n_2316;
     end
 assign n_1016 = retime_s9_35_reg_reg_IQ;
 reg retime_s9_37_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_37_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_37_reg_reg_IQ <= n_698;
     end
 assign n_697 = retime_s9_37_reg_reg_IQ;
 reg retime_s9_38_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_38_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_38_reg_reg_IQ <= n_686;
     end
 assign n_685 = retime_s9_38_reg_reg_IQ;
 reg retime_s9_39_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_39_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_39_reg_reg_IQ <= n_676;
     end
 assign n_675 = retime_s9_39_reg_reg_IQ;
 reg retime_s9_40_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_40_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_40_reg_reg_IQ <= n_169;
     end
 assign n_673 = retime_s9_40_reg_reg_IQ;
 reg retime_s9_41_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_41_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_41_reg_reg_IQ <= n_663;
     end
 assign n_662 = retime_s9_41_reg_reg_IQ;
 reg retime_s9_42_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_42_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_42_reg_reg_IQ <= n_653;
     end
 assign n_652 = retime_s9_42_reg_reg_IQ;
 reg retime_s9_43_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_43_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_43_reg_reg_IQ <= n_635;
     end
 assign n_634 = retime_s9_43_reg_reg_IQ;
 reg retime_s9_44_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_44_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_44_reg_reg_IQ <= n_621;
     end
 assign n_620 = retime_s9_44_reg_reg_IQ;
 reg retime_s9_45_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_45_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_45_reg_reg_IQ <= n_607;
     end
 assign n_606 = retime_s9_45_reg_reg_IQ;
 reg retime_s9_46_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_46_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_46_reg_reg_IQ <= n_597;
     end
 assign n_596 = retime_s9_46_reg_reg_IQ;
 reg retime_s9_47_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_47_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_47_reg_reg_IQ <= n_587;
     end
 assign n_586 = retime_s9_47_reg_reg_IQ;
 reg retime_s9_48_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_48_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_48_reg_reg_IQ <= n_561;
     end
 assign n_560 = retime_s9_48_reg_reg_IQ;
 reg retime_s9_49_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_49_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_49_reg_reg_IQ <= n_551;
     end
 assign n_550 = retime_s9_49_reg_reg_IQ;
 reg retime_s9_50_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_50_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_50_reg_reg_IQ <= n_541;
     end
 assign n_540 = retime_s9_50_reg_reg_IQ;
 reg retime_s9_51_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_51_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_51_reg_reg_IQ <= n_531;
     end
 assign n_530 = retime_s9_51_reg_reg_IQ;
 reg retime_s9_52_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_52_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_52_reg_reg_IQ <= n_520;
     end
 assign n_519 = retime_s9_52_reg_reg_IQ;
 reg retime_s9_53_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_53_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_53_reg_reg_IQ <= n_170;
     end
 assign n_511 = retime_s9_53_reg_reg_IQ;
 reg retime_s9_55_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_55_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_55_reg_reg_IQ <= n_114;
     end
 assign n_509 = retime_s9_55_reg_reg_IQ;
 reg retime_s9_56_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_56_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_56_reg_reg_IQ <= n_275;
     end
 assign n_508 = retime_s9_56_reg_reg_IQ;
 reg retime_s9_57_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_57_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_57_reg_reg_IQ <= n_500;
     end
 assign n_499 = retime_s9_57_reg_reg_IQ;
 reg retime_s9_58_reg_reg_IQ;
 wire retime_s9_58_reg_reg_IQN;
 assign retime_s9_58_reg_reg_IQN = !retime_s9_58_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_58_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_58_reg_reg_IQ <= n_162;
     end
 assign n_274 = retime_s9_58_reg_reg_IQN;
 reg retime_s9_59_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_59_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_59_reg_reg_IQ <= n_479;
     end
 assign n_478 = retime_s9_59_reg_reg_IQ;
 reg retime_s9_60_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_60_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_60_reg_reg_IQ <= n_469;
     end
 assign n_468 = retime_s9_60_reg_reg_IQ;
 reg retime_s9_61_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_61_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_61_reg_reg_IQ <= n_459;
     end
 assign n_458 = retime_s9_61_reg_reg_IQ;
 reg retime_s9_62_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_62_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_62_reg_reg_IQ <= n_449;
     end
 assign n_448 = retime_s9_62_reg_reg_IQ;
 reg retime_s9_63_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_63_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_63_reg_reg_IQ <= n_438;
     end
 assign n_437 = retime_s9_63_reg_reg_IQ;
 reg retime_s9_64_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_64_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_64_reg_reg_IQ <= n_428;
     end
 assign n_427 = retime_s9_64_reg_reg_IQ;
 reg retime_s9_65_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_65_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_65_reg_reg_IQ <= n_418;
     end
 assign n_417 = retime_s9_65_reg_reg_IQ;
 reg retime_s9_66_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_66_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_66_reg_reg_IQ <= n_408;
     end
 assign n_407 = retime_s9_66_reg_reg_IQ;
 reg retime_s9_67_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_67_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_67_reg_reg_IQ <= n_394;
     end
 assign n_393 = retime_s9_67_reg_reg_IQ;
 reg retime_s9_68_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_68_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_68_reg_reg_IQ <= n_384;
     end
 assign n_383 = retime_s9_68_reg_reg_IQ;
 reg retime_s9_69_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_69_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_69_reg_reg_IQ <= n_369;
     end
 assign n_368 = retime_s9_69_reg_reg_IQ;
 reg retime_s9_70_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_70_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_70_reg_reg_IQ <= n_358;
     end
 assign n_357 = retime_s9_70_reg_reg_IQ;
 reg retime_s9_71_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_71_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_71_reg_reg_IQ <= n_348;
     end
 assign n_347 = retime_s9_71_reg_reg_IQ;
 reg retime_s9_72_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_72_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_72_reg_reg_IQ <= n_337;
     end
 assign n_336 = retime_s9_72_reg_reg_IQ;
 reg retime_s10_1_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_1_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_1_reg_reg_IQ <= n_176;
     end
 assign n_1117 = retime_s10_1_reg_reg_IQ;
 reg retime_s10_2_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_2_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_2_reg_reg_IQ <= n_159;
     end
 assign n_1116 = retime_s10_2_reg_reg_IQ;
 reg retime_s10_3_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_3_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_3_reg_reg_IQ <= n_1107;
     end
 assign n_1106 = retime_s10_3_reg_reg_IQ;
 reg retime_s10_4_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_4_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_4_reg_reg_IQ <= n_2375;
     end
 assign n_1105 = retime_s10_4_reg_reg_IQ;
 reg retime_s10_5_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_5_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_5_reg_reg_IQ <= n_2383;
     end
 assign n_1104 = retime_s10_5_reg_reg_IQ;
 reg retime_s10_6_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_6_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_6_reg_reg_IQ <= n_2395;
     end
 assign n_1103 = retime_s10_6_reg_reg_IQ;
 reg retime_s10_7_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_7_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_7_reg_reg_IQ <= n_2396;
     end
 assign n_1102 = retime_s10_7_reg_reg_IQ;
 reg retime_s10_8_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_8_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_8_reg_reg_IQ <= sub_732_2_n_14;
     end
 assign n_1101 = retime_s10_8_reg_reg_IQ;
 reg retime_s10_9_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_9_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_9_reg_reg_IQ <= n_2427;
     end
 assign n_1100 = retime_s10_9_reg_reg_IQ;
 reg retime_s10_10_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_10_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_10_reg_reg_IQ <= n_2426;
     end
 assign n_1099 = retime_s10_10_reg_reg_IQ;
 reg retime_s10_11_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_11_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_11_reg_reg_IQ <= n_2425;
     end
 assign n_1098 = retime_s10_11_reg_reg_IQ;
 reg retime_s10_12_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_12_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_12_reg_reg_IQ <= n_2424;
     end
 assign n_1097 = retime_s10_12_reg_reg_IQ;
 reg retime_s10_13_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_13_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_13_reg_reg_IQ <= sub_732_2_n_156;
     end
 assign n_1096 = retime_s10_13_reg_reg_IQ;
 reg retime_s10_14_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_14_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_14_reg_reg_IQ <= n_2422;
     end
 assign n_1095 = retime_s10_14_reg_reg_IQ;
 reg retime_s10_15_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_15_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_15_reg_reg_IQ <= n_2423;
     end
 assign n_1094 = retime_s10_15_reg_reg_IQ;
 reg retime_s10_16_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_16_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_16_reg_reg_IQ <= n_2420;
     end
 assign n_1093 = retime_s10_16_reg_reg_IQ;
 reg retime_s10_17_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_17_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_17_reg_reg_IQ <= n_2419;
     end
 assign n_1092 = retime_s10_17_reg_reg_IQ;
 reg retime_s10_18_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_18_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_18_reg_reg_IQ <= sub_732_2_n_172;
     end
 assign n_1091 = retime_s10_18_reg_reg_IQ;
 reg retime_s10_19_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_19_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_19_reg_reg_IQ <= n_2418;
     end
 assign n_1090 = retime_s10_19_reg_reg_IQ;
 reg retime_s10_20_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_20_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_20_reg_reg_IQ <= n_2421;
     end
 assign n_1089 = retime_s10_20_reg_reg_IQ;
 reg retime_s10_21_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_21_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_21_reg_reg_IQ <= n_2394;
     end
 assign n_1088 = retime_s10_21_reg_reg_IQ;
 reg retime_s10_22_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_22_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_22_reg_reg_IQ <= n_2374;
     end
 assign n_1087 = retime_s10_22_reg_reg_IQ;
 reg retime_s10_23_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_23_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_23_reg_reg_IQ <= n_2393;
     end
 assign n_1086 = retime_s10_23_reg_reg_IQ;
 reg retime_s10_24_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_24_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_24_reg_reg_IQ <= n_2380;
     end
 assign n_1085 = retime_s10_24_reg_reg_IQ;
 reg retime_s10_25_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_25_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_25_reg_reg_IQ <= n_2376;
     end
 assign n_1084 = retime_s10_25_reg_reg_IQ;
 reg retime_s10_26_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_26_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_26_reg_reg_IQ <= n_2390;
     end
 assign n_1083 = retime_s10_26_reg_reg_IQ;
 reg retime_s10_27_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_27_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_27_reg_reg_IQ <= sub_732_2_n_54;
     end
 assign n_1082 = retime_s10_27_reg_reg_IQ;
 reg retime_s10_28_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_28_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_28_reg_reg_IQ <= n_2373;
     end
 assign n_1081 = retime_s10_28_reg_reg_IQ;
 reg retime_s10_29_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_29_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_29_reg_reg_IQ <= n_2391;
     end
 assign n_1080 = retime_s10_29_reg_reg_IQ;
 reg retime_s10_30_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_30_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_30_reg_reg_IQ <= n_2400;
     end
 assign n_1079 = retime_s10_30_reg_reg_IQ;
 reg retime_s10_31_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_31_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_31_reg_reg_IQ <= n_2431;
     end
 assign n_1078 = retime_s10_31_reg_reg_IQ;
 reg retime_s10_32_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_32_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_32_reg_reg_IQ <= n_2429;
     end
 assign n_1077 = retime_s10_32_reg_reg_IQ;
 reg retime_s10_33_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_33_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_33_reg_reg_IQ <= n_2428;
     end
 assign n_1076 = retime_s10_33_reg_reg_IQ;
 reg retime_s10_34_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_34_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_34_reg_reg_IQ <= n_2430;
     end
 assign n_1075 = retime_s10_34_reg_reg_IQ;
 reg retime_s10_35_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_35_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_35_reg_reg_IQ <= n_2378;
     end
 assign n_1074 = retime_s10_35_reg_reg_IQ;
 reg retime_s10_36_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_36_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_36_reg_reg_IQ <= n_2372;
     end
 assign n_1073 = retime_s10_36_reg_reg_IQ;
 reg retime_s10_37_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_37_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_37_reg_reg_IQ <= n_2389;
     end
 assign n_1072 = retime_s10_37_reg_reg_IQ;
 reg retime_s10_38_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_38_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_38_reg_reg_IQ <= n_2397;
     end
 assign n_1071 = retime_s10_38_reg_reg_IQ;
 reg retime_s10_39_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_39_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_39_reg_reg_IQ <= n_2398;
     end
 assign n_1070 = retime_s10_39_reg_reg_IQ;
 reg retime_s10_40_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_40_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_40_reg_reg_IQ <= n_2399;
     end
 assign n_1069 = retime_s10_40_reg_reg_IQ;
 reg retime_s10_41_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_41_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_41_reg_reg_IQ <= n_2371;
     end
 assign n_1068 = retime_s10_41_reg_reg_IQ;
 reg retime_s10_42_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_42_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_42_reg_reg_IQ <= n_2387;
     end
 assign n_1067 = retime_s10_42_reg_reg_IQ;
 reg retime_s10_43_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_43_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_43_reg_reg_IQ <= n_2379;
     end
 assign n_1066 = retime_s10_43_reg_reg_IQ;
 reg retime_s10_44_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_44_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_44_reg_reg_IQ <= sub_732_2_n_16;
     end
 assign n_1065 = retime_s10_44_reg_reg_IQ;
 reg retime_s10_45_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_45_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_45_reg_reg_IQ <= n_2385;
     end
 assign n_1064 = retime_s10_45_reg_reg_IQ;
 reg retime_s10_46_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_46_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_46_reg_reg_IQ <= n_2377;
     end
 assign n_1063 = retime_s10_46_reg_reg_IQ;
 reg retime_s10_47_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_47_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_47_reg_reg_IQ <= sub_732_2_n_34;
     end
 assign n_1062 = retime_s10_47_reg_reg_IQ;
 reg retime_s10_48_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_48_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_48_reg_reg_IQ <= sub_732_2_n_36;
     end
 assign n_1061 = retime_s10_48_reg_reg_IQ;
 reg retime_s10_49_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_49_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_49_reg_reg_IQ <= n_2386;
     end
 assign n_1060 = retime_s10_49_reg_reg_IQ;
 reg retime_s10_50_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_50_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_50_reg_reg_IQ <= n_2381;
     end
 assign n_1059 = retime_s10_50_reg_reg_IQ;
 reg retime_s10_51_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_51_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_51_reg_reg_IQ <= n_2388;
     end
 assign n_1058 = retime_s10_51_reg_reg_IQ;
 reg retime_s10_52_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_52_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_52_reg_reg_IQ <= sub_732_2_n_11;
     end
 assign n_1057 = retime_s10_52_reg_reg_IQ;
 reg retime_s10_53_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_53_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_53_reg_reg_IQ <= sub_732_2_n_35;
     end
 assign n_1056 = retime_s10_53_reg_reg_IQ;
 reg retime_s10_54_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_54_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_54_reg_reg_IQ <= sub_732_2_n_91;
     end
 assign n_1055 = retime_s10_54_reg_reg_IQ;
 reg retime_s10_55_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_55_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_55_reg_reg_IQ <= sub_732_2_n_8;
     end
 assign n_1054 = retime_s10_55_reg_reg_IQ;
 reg retime_s10_56_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_56_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_56_reg_reg_IQ <= n_2384;
     end
 assign n_1053 = retime_s10_56_reg_reg_IQ;
 reg retime_s10_57_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_57_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_57_reg_reg_IQ <= n_2382;
     end
 assign n_1052 = retime_s10_57_reg_reg_IQ;
 reg retime_s10_58_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_58_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_58_reg_reg_IQ <= sub_732_2_n_25;
     end
 assign n_1051 = retime_s10_58_reg_reg_IQ;
 reg retime_s10_59_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_59_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_59_reg_reg_IQ <= sub_732_2_n_21;
     end
 assign n_1050 = retime_s10_59_reg_reg_IQ;
 reg retime_s10_60_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_60_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_60_reg_reg_IQ <= sub_732_2_n_6;
     end
 assign n_1049 = retime_s10_60_reg_reg_IQ;
 reg retime_s10_61_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_61_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_61_reg_reg_IQ <= n_2392;
     end
 assign n_1048 = retime_s10_61_reg_reg_IQ;
 reg retime_s10_62_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_62_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_62_reg_reg_IQ <= n_223;
     end
 assign n_706 = retime_s10_62_reg_reg_IQ;
 reg retime_s10_63_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_63_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_63_reg_reg_IQ <= n_697;
     end
 assign n_696 = retime_s10_63_reg_reg_IQ;
 reg retime_s10_64_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_64_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_64_reg_reg_IQ <= n_685;
     end
 assign n_684 = retime_s10_64_reg_reg_IQ;
 reg retime_s10_65_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_65_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_65_reg_reg_IQ <= n_675;
     end
 assign n_674 = retime_s10_65_reg_reg_IQ;
 reg retime_s10_66_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_66_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_66_reg_reg_IQ <= n_662;
     end
 assign n_661 = retime_s10_66_reg_reg_IQ;
 reg retime_s10_67_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_67_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_67_reg_reg_IQ <= n_652;
     end
 assign n_651 = retime_s10_67_reg_reg_IQ;
 reg retime_s10_68_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_68_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_68_reg_reg_IQ <= n_634;
     end
 assign n_633 = retime_s10_68_reg_reg_IQ;
 reg retime_s10_69_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_69_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_69_reg_reg_IQ <= n_620;
     end
 assign n_619 = retime_s10_69_reg_reg_IQ;
 reg retime_s10_70_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_70_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_70_reg_reg_IQ <= n_606;
     end
 assign n_605 = retime_s10_70_reg_reg_IQ;
 reg retime_s10_71_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_71_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_71_reg_reg_IQ <= n_596;
     end
 assign n_595 = retime_s10_71_reg_reg_IQ;
 reg retime_s10_72_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_72_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_72_reg_reg_IQ <= n_586;
     end
 assign n_585 = retime_s10_72_reg_reg_IQ;
 reg retime_s10_73_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_73_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_73_reg_reg_IQ <= n_560;
     end
 assign n_559 = retime_s10_73_reg_reg_IQ;
 reg retime_s10_74_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_74_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_74_reg_reg_IQ <= n_550;
     end
 assign n_549 = retime_s10_74_reg_reg_IQ;
 reg retime_s10_75_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_75_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_75_reg_reg_IQ <= n_540;
     end
 assign n_539 = retime_s10_75_reg_reg_IQ;
 reg retime_s10_76_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_76_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_76_reg_reg_IQ <= n_530;
     end
 assign n_529 = retime_s10_76_reg_reg_IQ;
 reg retime_s10_77_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_77_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_77_reg_reg_IQ <= n_519;
     end
 assign n_518 = retime_s10_77_reg_reg_IQ;
 reg retime_s10_78_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_78_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_78_reg_reg_IQ <= n_105;
     end
 assign n_510 = retime_s10_78_reg_reg_IQ;
 reg retime_s10_79_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_79_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_79_reg_reg_IQ <= n_499;
     end
 assign n_498 = retime_s10_79_reg_reg_IQ;
 reg retime_s10_80_reg_reg_IQ;
 wire retime_s10_80_reg_reg_IQN;
 assign retime_s10_80_reg_reg_IQN = !retime_s10_80_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_80_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_80_reg_reg_IQ <= n_274;
     end
 assign n_497 = retime_s10_80_reg_reg_IQN;
 reg retime_s10_81_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_81_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_81_reg_reg_IQ <= n_478;
     end
 assign n_477 = retime_s10_81_reg_reg_IQ;
 reg retime_s10_82_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_82_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_82_reg_reg_IQ <= n_468;
     end
 assign n_467 = retime_s10_82_reg_reg_IQ;
 reg retime_s10_83_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_83_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_83_reg_reg_IQ <= n_458;
     end
 assign n_457 = retime_s10_83_reg_reg_IQ;
 reg retime_s10_84_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_84_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_84_reg_reg_IQ <= n_448;
     end
 assign n_447 = retime_s10_84_reg_reg_IQ;
 reg retime_s10_85_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_85_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_85_reg_reg_IQ <= n_437;
     end
 assign n_436 = retime_s10_85_reg_reg_IQ;
 reg retime_s10_86_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_86_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_86_reg_reg_IQ <= n_427;
     end
 assign n_426 = retime_s10_86_reg_reg_IQ;
 reg retime_s10_87_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_87_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_87_reg_reg_IQ <= n_417;
     end
 assign n_416 = retime_s10_87_reg_reg_IQ;
 reg retime_s10_88_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_88_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_88_reg_reg_IQ <= n_407;
     end
 assign n_406 = retime_s10_88_reg_reg_IQ;
 reg retime_s10_89_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_89_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_89_reg_reg_IQ <= n_393;
     end
 assign n_392 = retime_s10_89_reg_reg_IQ;
 reg retime_s10_90_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_90_reg_reg_IQ <= 1'B0;
     else begin
         retime_s10_90_reg_reg_IQ <= sub_751_2_n_0;
     end
 assign n_382 = retime_s10_90_reg_reg_IQ;
 reg retime_s10_91_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_91_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_91_reg_reg_IQ <= n_368;
     end
 assign n_367 = retime_s10_91_reg_reg_IQ;
 reg retime_s10_92_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_92_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_92_reg_reg_IQ <= n_357;
     end
 assign n_356 = retime_s10_92_reg_reg_IQ;
 reg retime_s10_93_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_93_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_93_reg_reg_IQ <= n_347;
     end
 assign n_346 = retime_s10_93_reg_reg_IQ;
 reg retime_s10_94_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s10_94_reg_reg_IQ <= 1'B1;
     else begin
         retime_s10_94_reg_reg_IQ <= n_336;
     end
 assign n_335 = retime_s10_94_reg_reg_IQ;
 reg retime_s1_1_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_1_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_1_reg_reg_IQ <= {in2[0]};
     end
 assign n_156 = retime_s1_1_reg_reg_IQ;
 reg retime_s1_2_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_2_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_2_reg_reg_IQ <= {in2[1]};
     end
 assign n_182 = retime_s1_2_reg_reg_IQ;
 reg retime_s1_7_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_7_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_7_reg_reg_IQ <= {in2[21]};
     end
 assign n_155 = retime_s1_7_reg_reg_IQ;
 reg retime_s1_8_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_8_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_8_reg_reg_IQ <= n_1572;
     end
 assign n_101 = retime_s1_8_reg_reg_IQ;
 reg retime_s1_10_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_10_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_10_reg_reg_IQ <= {in2[6]};
     end
 assign n_154 = retime_s1_10_reg_reg_IQ;
 reg retime_s1_11_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_11_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_11_reg_reg_IQ <= sub_637_2_n_35;
     end
 assign n_102 = retime_s1_11_reg_reg_IQ;
 reg retime_s1_13_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_13_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_13_reg_reg_IQ <= {in2[16]};
     end
 assign n_85 = retime_s1_13_reg_reg_IQ;
 reg retime_s1_14_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_14_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_14_reg_reg_IQ <= sub_352_2_n_36;
     end
 assign n_153 = retime_s1_14_reg_reg_IQ;
 reg retime_s1_15_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_15_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_15_reg_reg_IQ <= sub_447_2_n_56;
     end
 assign n_76 = retime_s1_15_reg_reg_IQ;
 reg retime_s1_16_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_16_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_16_reg_reg_IQ <= n_1712;
     end
 assign n_152 = retime_s1_16_reg_reg_IQ;
 reg retime_s1_20_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_20_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_20_reg_reg_IQ <= {in2[10]};
     end
 assign n_96 = retime_s1_20_reg_reg_IQ;
 reg retime_s1_21_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_21_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_21_reg_reg_IQ <= sub_561_2_n_55;
     end
 assign n_80 = retime_s1_21_reg_reg_IQ;
 reg retime_s1_24_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_24_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_24_reg_reg_IQ <= n_2432;
     end
 assign n_150 = retime_s1_24_reg_reg_IQ;
 reg retime_s1_30_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_30_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_30_reg_reg_IQ <= sub_732_2_n_33;
     end
 assign n_86 = retime_s1_30_reg_reg_IQ;
 reg retime_s1_31_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_31_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_31_reg_reg_IQ <= n_1946;
     end
 assign n_178 = retime_s1_31_reg_reg_IQ;
 reg retime_s1_32_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_32_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_32_reg_reg_IQ <= {in2[13]};
     end
 assign n_179 = retime_s1_32_reg_reg_IQ;
 reg retime_s1_35_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_35_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_35_reg_reg_IQ <= n_1820;
     end
 assign n_181 = retime_s1_35_reg_reg_IQ;
 reg retime_s1_44_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_44_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_44_reg_reg_IQ <= {in2[18]};
     end
 assign n_183 = retime_s1_44_reg_reg_IQ;
 reg retime_s1_45_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_45_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_45_reg_reg_IQ <= sub_409_2_n_35;
     end
 assign n_184 = retime_s1_45_reg_reg_IQ;
 reg retime_s1_46_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_46_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_46_reg_reg_IQ <= n_1650;
     end
 assign n_185 = retime_s1_46_reg_reg_IQ;
 reg retime_s1_47_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_47_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_47_reg_reg_IQ <= {in2[12]};
     end
 assign n_186 = retime_s1_47_reg_reg_IQ;
 reg retime_s1_49_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_49_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_49_reg_reg_IQ <= {in2[17]};
     end
 assign n_187 = retime_s1_49_reg_reg_IQ;
 reg retime_s1_51_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_51_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_51_reg_reg_IQ <= sub_428_2_n_54;
     end
 assign n_188 = retime_s1_51_reg_reg_IQ;
 reg retime_s1_52_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_52_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_52_reg_reg_IQ <= n_1680;
     end
 assign n_190 = retime_s1_52_reg_reg_IQ;
 reg retime_s1_56_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_56_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_56_reg_reg_IQ <= {in2[19]};
     end
 assign n_191 = retime_s1_56_reg_reg_IQ;
 reg retime_s1_57_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_57_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_57_reg_reg_IQ <= sub_390_2_n_45;
     end
 assign n_192 = retime_s1_57_reg_reg_IQ;
 reg retime_s1_58_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_58_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_58_reg_reg_IQ <= n_1622;
     end
 assign n_193 = retime_s1_58_reg_reg_IQ;
 reg retime_s1_59_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_59_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_59_reg_reg_IQ <= {in2[20]};
     end
 assign n_194 = retime_s1_59_reg_reg_IQ;
 reg retime_s1_60_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_60_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_60_reg_reg_IQ <= n_1596;
     end
 assign n_195 = retime_s1_60_reg_reg_IQ;
 reg retime_s1_61_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_61_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_61_reg_reg_IQ <= sub_371_2_n_26;
     end
 assign n_196 = retime_s1_61_reg_reg_IQ;
 reg retime_s1_62_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_62_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_62_reg_reg_IQ <= {in2[22]};
     end
 assign n_197 = retime_s1_62_reg_reg_IQ;
 reg retime_s1_65_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_65_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_65_reg_reg_IQ <= n_1860;
     end
 assign n_198 = retime_s1_65_reg_reg_IQ;
 reg retime_s1_66_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_66_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_66_reg_reg_IQ <= {in2[9]};
     end
 assign n_199 = retime_s1_66_reg_reg_IQ;
 reg retime_s1_67_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_67_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_67_reg_reg_IQ <= {in2[5]};
     end
 assign n_200 = retime_s1_67_reg_reg_IQ;
 reg retime_s1_68_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_68_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_68_reg_reg_IQ <= sub_580_2_n_59;
     end
 assign n_201 = retime_s1_68_reg_reg_IQ;
 reg retime_s1_69_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_69_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_69_reg_reg_IQ <= sub_656_2_n_64;
     end
 assign n_202 = retime_s1_69_reg_reg_IQ;
 reg retime_s1_70_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_70_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_70_reg_reg_IQ <= n_2196;
     end
 assign n_203 = retime_s1_70_reg_reg_IQ;
 reg retime_s1_71_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_71_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_71_reg_reg_IQ <= n_1992;
     end
 assign n_204 = retime_s1_71_reg_reg_IQ;
 reg retime_s1_78_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_78_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_78_reg_reg_IQ <= {in2[3]};
     end
 assign n_206 = retime_s1_78_reg_reg_IQ;
 reg retime_s1_79_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_79_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_79_reg_reg_IQ <= sub_694_2_n_39;
     end
 assign n_207 = retime_s1_79_reg_reg_IQ;
 reg retime_s1_80_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_80_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_80_reg_reg_IQ <= n_2310;
     end
 assign n_208 = retime_s1_80_reg_reg_IQ;
 reg retime_s1_81_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_81_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_81_reg_reg_IQ <= {in2[8]};
     end
 assign n_209 = retime_s1_81_reg_reg_IQ;
 reg retime_s1_82_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_82_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_82_reg_reg_IQ <= sub_599_2_n_48;
     end
 assign n_210 = retime_s1_82_reg_reg_IQ;
 reg retime_s1_83_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_83_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_83_reg_reg_IQ <= n_2040;
     end
 assign n_211 = retime_s1_83_reg_reg_IQ;
 reg retime_s1_84_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_84_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_84_reg_reg_IQ <= {in2[2]};
     end
 assign n_212 = retime_s1_84_reg_reg_IQ;
 reg retime_s1_85_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_85_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_85_reg_reg_IQ <= n_2496;
     end
 assign n_213 = retime_s1_85_reg_reg_IQ;
 reg retime_s1_86_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_86_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_86_reg_reg_IQ <= sub_713_2_n_4;
     end
 assign n_214 = retime_s1_86_reg_reg_IQ;
 reg retime_s1_87_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_87_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_87_reg_reg_IQ <= n_2370;
     end
 assign n_215 = retime_s1_87_reg_reg_IQ;
 reg retime_s1_89_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_89_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_89_reg_reg_IQ <= sub_751_2_n_1;
     end
 assign n_216 = retime_s1_89_reg_reg_IQ;
 reg retime_s1_90_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_90_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_90_reg_reg_IQ <= {in2[11]};
     end
 assign n_217 = retime_s1_90_reg_reg_IQ;
 reg retime_s1_91_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_91_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_91_reg_reg_IQ <= sub_542_2_n_52;
     end
 assign n_218 = retime_s1_91_reg_reg_IQ;
 reg retime_s1_93_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_93_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_93_reg_reg_IQ <= n_1902;
     end
 assign n_219 = retime_s1_93_reg_reg_IQ;
 reg retime_s1_94_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_94_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_94_reg_reg_IQ <= {in2[15]};
     end
 assign n_220 = retime_s1_94_reg_reg_IQ;
 reg retime_s1_95_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_95_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_95_reg_reg_IQ <= sub_466_2_n_52;
     end
 assign n_221 = retime_s1_95_reg_reg_IQ;
 reg retime_s1_96_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_96_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_96_reg_reg_IQ <= n_1746;
     end
 assign n_222 = retime_s1_96_reg_reg_IQ;
 reg retime_s1_104_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_104_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_104_reg_reg_IQ <= n_2142;
     end
 assign n_224 = retime_s1_104_reg_reg_IQ;
 reg retime_s1_109_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_109_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_109_reg_reg_IQ <= {in2[14]};
     end
 assign n_225 = retime_s1_109_reg_reg_IQ;
 reg retime_s1_110_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_110_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_110_reg_reg_IQ <= sub_485_2_n_32;
     end
 assign n_226 = retime_s1_110_reg_reg_IQ;
 reg retime_s1_111_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_111_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_111_reg_reg_IQ <= n_1782;
     end
 assign n_227 = retime_s1_111_reg_reg_IQ;
 reg retime_s1_112_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_112_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_112_reg_reg_IQ <= sub_523_2_n_52;
     end
 assign n_228 = retime_s1_112_reg_reg_IQ;
 reg retime_s1_115_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_115_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_115_reg_reg_IQ <= sub_504_2_n_29;
     end
 assign n_229 = retime_s1_115_reg_reg_IQ;
 reg retime_s1_116_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_116_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_116_reg_reg_IQ <= sub_675_2_n_29;
     end
 assign n_230 = retime_s1_116_reg_reg_IQ;
 reg retime_s1_117_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_117_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_117_reg_reg_IQ <= n_2252;
     end
 assign n_231 = retime_s1_117_reg_reg_IQ;
 reg retime_s1_118_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_118_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_118_reg_reg_IQ <= sub_618_2_n_48;
     end
 assign n_232 = retime_s1_118_reg_reg_IQ;
 reg retime_s1_119_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_119_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_119_reg_reg_IQ <= n_2090;
     end
 assign n_233 = retime_s1_119_reg_reg_IQ;
 reg retime_s1_121_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_121_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_121_reg_reg_IQ <= {in2[4]};
     end
 assign n_234 = retime_s1_121_reg_reg_IQ;
 reg retime_s1_124_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_124_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_124_reg_reg_IQ <= {in2[7]};
     end
 assign n_235 = retime_s1_124_reg_reg_IQ;
 reg retime_s2_1_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_1_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_1_reg_reg_IQ <= n_156;
     end
 assign n_236 = retime_s2_1_reg_reg_IQ;
 reg retime_s2_2_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_2_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_2_reg_reg_IQ <= n_182;
     end
 assign n_237 = retime_s2_2_reg_reg_IQ;
 reg retime_s2_30_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_30_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_30_reg_reg_IQ <= n_154;
     end
 assign n_239 = retime_s2_30_reg_reg_IQ;
 reg retime_s2_31_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_31_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_31_reg_reg_IQ <= n_102;
     end
 assign n_240 = retime_s2_31_reg_reg_IQ;
 reg retime_s2_32_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_32_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_32_reg_reg_IQ <= n_85;
     end
 assign n_241 = retime_s2_32_reg_reg_IQ;
 reg retime_s2_34_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_34_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_34_reg_reg_IQ <= n_76;
     end
 assign n_242 = retime_s2_34_reg_reg_IQ;
 reg retime_s2_35_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_35_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_35_reg_reg_IQ <= n_152;
     end
 assign n_243 = retime_s2_35_reg_reg_IQ;
 reg retime_s2_36_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_36_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_36_reg_reg_IQ <= n_96;
     end
 assign n_244 = retime_s2_36_reg_reg_IQ;
 reg retime_s2_37_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_37_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_37_reg_reg_IQ <= n_80;
     end
 assign n_245 = retime_s2_37_reg_reg_IQ;
 reg retime_s2_38_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_38_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_38_reg_reg_IQ <= n_150;
     end
 assign n_246 = retime_s2_38_reg_reg_IQ;
 reg retime_s2_42_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_42_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_42_reg_reg_IQ <= n_86;
     end
 assign n_248 = retime_s2_42_reg_reg_IQ;
 reg retime_s2_43_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_43_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_43_reg_reg_IQ <= n_178;
     end
 assign n_249 = retime_s2_43_reg_reg_IQ;
 reg retime_s2_44_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_44_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_44_reg_reg_IQ <= n_179;
     end
 assign n_250 = retime_s2_44_reg_reg_IQ;
 reg retime_s2_47_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_47_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_47_reg_reg_IQ <= n_181;
     end
 assign n_251 = retime_s2_47_reg_reg_IQ;
 reg retime_s2_49_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_49_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_49_reg_reg_IQ <= n_183;
     end
 assign n_252 = retime_s2_49_reg_reg_IQ;
 reg retime_s2_50_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_50_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_50_reg_reg_IQ <= n_184;
     end
 assign n_253 = retime_s2_50_reg_reg_IQ;
 reg retime_s2_51_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_51_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_51_reg_reg_IQ <= n_185;
     end
 assign n_254 = retime_s2_51_reg_reg_IQ;
 reg retime_s2_52_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_52_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_52_reg_reg_IQ <= n_186;
     end
 assign n_255 = retime_s2_52_reg_reg_IQ;
 reg retime_s2_54_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_54_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_54_reg_reg_IQ <= n_187;
     end
 assign n_256 = retime_s2_54_reg_reg_IQ;
 reg retime_s2_55_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_55_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_55_reg_reg_IQ <= n_188;
     end
 assign n_257 = retime_s2_55_reg_reg_IQ;
 reg retime_s2_56_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_56_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_56_reg_reg_IQ <= n_190;
     end
 assign n_258 = retime_s2_56_reg_reg_IQ;
 reg retime_s2_60_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_60_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_60_reg_reg_IQ <= n_191;
     end
 assign n_259 = retime_s2_60_reg_reg_IQ;
 reg retime_s2_62_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_62_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_62_reg_reg_IQ <= n_193;
     end
 assign n_260 = retime_s2_62_reg_reg_IQ;
 reg retime_s2_68_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_68_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_68_reg_reg_IQ <= n_198;
     end
 assign n_261 = retime_s2_68_reg_reg_IQ;
 reg retime_s2_69_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_69_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_69_reg_reg_IQ <= n_199;
     end
 assign n_262 = retime_s2_69_reg_reg_IQ;
 reg retime_s2_70_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_70_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_70_reg_reg_IQ <= n_200;
     end
 assign n_263 = retime_s2_70_reg_reg_IQ;
 reg retime_s2_71_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_71_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_71_reg_reg_IQ <= n_201;
     end
 assign n_264 = retime_s2_71_reg_reg_IQ;
 reg retime_s2_72_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_72_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_72_reg_reg_IQ <= n_202;
     end
 assign n_265 = retime_s2_72_reg_reg_IQ;
 reg retime_s2_73_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_73_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_73_reg_reg_IQ <= n_203;
     end
 assign n_266 = retime_s2_73_reg_reg_IQ;
 reg retime_s2_74_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_74_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_74_reg_reg_IQ <= n_204;
     end
 assign n_267 = retime_s2_74_reg_reg_IQ;
 reg retime_s2_80_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_80_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_80_reg_reg_IQ <= n_206;
     end
 assign n_136 = retime_s2_80_reg_reg_IQ;
 reg retime_s2_81_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_81_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_81_reg_reg_IQ <= n_207;
     end
 assign n_130 = retime_s2_81_reg_reg_IQ;
 reg retime_s2_82_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_82_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_82_reg_reg_IQ <= n_208;
     end
 assign n_87 = retime_s2_82_reg_reg_IQ;
 reg retime_s2_83_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_83_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_83_reg_reg_IQ <= n_209;
     end
 assign n_33 = retime_s2_83_reg_reg_IQ;
 reg retime_s2_84_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_84_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_84_reg_reg_IQ <= n_210;
     end
 assign n_144 = retime_s2_84_reg_reg_IQ;
 reg retime_s2_85_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_85_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_85_reg_reg_IQ <= n_211;
     end
 assign n_84 = retime_s2_85_reg_reg_IQ;
 reg retime_s2_86_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_86_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_86_reg_reg_IQ <= n_212;
     end
 assign n_88 = retime_s2_86_reg_reg_IQ;
 reg retime_s2_87_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_87_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_87_reg_reg_IQ <= n_213;
     end
 assign n_32 = retime_s2_87_reg_reg_IQ;
 reg retime_s2_88_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_88_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_88_reg_reg_IQ <= n_214;
     end
 assign n_1 = retime_s2_88_reg_reg_IQ;
 reg retime_s2_89_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_89_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_89_reg_reg_IQ <= n_215;
     end
 assign n_82 = retime_s2_89_reg_reg_IQ;
 reg retime_s2_91_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_91_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_91_reg_reg_IQ <= n_216;
     end
 assign n_92 = retime_s2_91_reg_reg_IQ;
 reg retime_s2_92_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_92_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_92_reg_reg_IQ <= n_217;
     end
 assign n_31 = retime_s2_92_reg_reg_IQ;
 reg retime_s2_93_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_93_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_93_reg_reg_IQ <= n_218;
     end
 assign n_140 = retime_s2_93_reg_reg_IQ;
 reg retime_s2_94_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_94_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_94_reg_reg_IQ <= n_219;
     end
 assign n_139 = retime_s2_94_reg_reg_IQ;
 reg retime_s2_95_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_95_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_95_reg_reg_IQ <= n_220;
     end
 assign n_79 = retime_s2_95_reg_reg_IQ;
 reg retime_s2_96_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_96_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_96_reg_reg_IQ <= n_221;
     end
 assign n_138 = retime_s2_96_reg_reg_IQ;
 reg retime_s2_97_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_97_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_97_reg_reg_IQ <= n_222;
     end
 assign n_0 = retime_s2_97_reg_reg_IQ;
 reg retime_s2_102_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_102_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_102_reg_reg_IQ <= n_224;
     end
 assign n_78 = retime_s2_102_reg_reg_IQ;
 reg retime_s2_107_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_107_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_107_reg_reg_IQ <= n_225;
     end
 assign n_99 = retime_s2_107_reg_reg_IQ;
 reg retime_s2_108_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_108_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_108_reg_reg_IQ <= n_226;
     end
 assign n_30 = retime_s2_108_reg_reg_IQ;
 reg retime_s2_109_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_109_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_109_reg_reg_IQ <= n_227;
     end
 assign n_137 = retime_s2_109_reg_reg_IQ;
 reg retime_s2_110_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_110_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_110_reg_reg_IQ <= n_228;
     end
 assign n_29 = retime_s2_110_reg_reg_IQ;
 reg retime_s2_113_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_113_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_113_reg_reg_IQ <= n_229;
     end
 assign n_77 = retime_s2_113_reg_reg_IQ;
 reg retime_s2_114_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_114_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_114_reg_reg_IQ <= n_230;
     end
 assign n_100 = retime_s2_114_reg_reg_IQ;
 reg retime_s2_115_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_115_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_115_reg_reg_IQ <= n_231;
     end
 assign n_28 = retime_s2_115_reg_reg_IQ;
 reg retime_s2_116_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_116_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_116_reg_reg_IQ <= n_232;
     end
 assign n_27 = retime_s2_116_reg_reg_IQ;
 reg retime_s2_117_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_117_reg_reg_IQ <= 1'B1;
     else begin
         retime_s2_117_reg_reg_IQ <= n_233;
     end
 assign n_26 = retime_s2_117_reg_reg_IQ;
 reg retime_s2_119_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_119_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_119_reg_reg_IQ <= n_234;
     end
 assign n_103 = retime_s2_119_reg_reg_IQ;
 reg retime_s2_122_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s2_122_reg_reg_IQ <= 1'B0;
     else begin
         retime_s2_122_reg_reg_IQ <= n_235;
     end
 assign n_148 = retime_s2_122_reg_reg_IQ;
 reg retime_s3_1_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_1_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_1_reg_reg_IQ <= n_236;
     end
 assign n_75 = retime_s3_1_reg_reg_IQ;
 reg retime_s3_2_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_2_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_2_reg_reg_IQ <= n_237;
     end
 assign n_25 = retime_s3_2_reg_reg_IQ;
 reg retime_s3_34_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_34_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_34_reg_reg_IQ <= n_239;
     end
 assign n_24 = retime_s3_34_reg_reg_IQ;
 reg retime_s3_35_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_35_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_35_reg_reg_IQ <= n_240;
     end
 assign n_171 = retime_s3_35_reg_reg_IQ;
 reg retime_s3_39_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_39_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_39_reg_reg_IQ <= n_244;
     end
 assign n_23 = retime_s3_39_reg_reg_IQ;
 reg retime_s3_40_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_40_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_40_reg_reg_IQ <= n_245;
     end
 assign n_174 = retime_s3_40_reg_reg_IQ;
 reg retime_s3_41_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_41_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_41_reg_reg_IQ <= n_246;
     end
 assign n_68 = retime_s3_41_reg_reg_IQ;
 reg retime_s3_45_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_45_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_45_reg_reg_IQ <= n_248;
     end
 assign n_67 = retime_s3_45_reg_reg_IQ;
 reg retime_s3_46_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_46_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_46_reg_reg_IQ <= n_249;
     end
 assign n_34 = retime_s3_46_reg_reg_IQ;
 reg retime_s3_47_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_47_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_47_reg_reg_IQ <= n_250;
     end
 assign n_66 = retime_s3_47_reg_reg_IQ;
 reg retime_s3_50_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_50_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_50_reg_reg_IQ <= n_251;
     end
 assign n_124 = retime_s3_50_reg_reg_IQ;
 reg retime_s3_55_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_55_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_55_reg_reg_IQ <= n_255;
     end
 assign n_22 = retime_s3_55_reg_reg_IQ;
 reg retime_s3_65_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_65_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_65_reg_reg_IQ <= n_261;
     end
 assign n_107 = retime_s3_65_reg_reg_IQ;
 reg retime_s3_66_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_66_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_66_reg_reg_IQ <= n_262;
     end
 assign n_20 = retime_s3_66_reg_reg_IQ;
 reg retime_s3_67_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_67_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_67_reg_reg_IQ <= n_263;
     end
 assign n_189 = retime_s3_67_reg_reg_IQ;
 reg retime_s3_68_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_68_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_68_reg_reg_IQ <= n_264;
     end
 assign n_40 = retime_s3_68_reg_reg_IQ;
 reg retime_s3_69_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_69_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_69_reg_reg_IQ <= n_265;
     end
 assign n_62 = retime_s3_69_reg_reg_IQ;
 reg retime_s3_70_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_70_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_70_reg_reg_IQ <= n_266;
     end
 assign n_112 = retime_s3_70_reg_reg_IQ;
 reg retime_s3_71_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_71_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_71_reg_reg_IQ <= n_267;
     end
 assign n_19 = retime_s3_71_reg_reg_IQ;
 reg retime_s3_77_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_77_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_77_reg_reg_IQ <= n_136;
     end
 assign n_115 = retime_s3_77_reg_reg_IQ;
 reg retime_s3_78_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_78_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_78_reg_reg_IQ <= n_130;
     end
 assign n_18 = retime_s3_78_reg_reg_IQ;
 reg retime_s3_79_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_79_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_79_reg_reg_IQ <= n_87;
     end
 assign n_61 = retime_s3_79_reg_reg_IQ;
 reg retime_s3_80_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_80_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_80_reg_reg_IQ <= n_33;
     end
 assign n_135 = retime_s3_80_reg_reg_IQ;
 reg retime_s3_81_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_81_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_81_reg_reg_IQ <= n_144;
     end
 assign n_125 = retime_s3_81_reg_reg_IQ;
 reg retime_s3_82_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_82_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_82_reg_reg_IQ <= n_84;
     end
 assign n_46 = retime_s3_82_reg_reg_IQ;
 reg retime_s3_83_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_83_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_83_reg_reg_IQ <= n_88;
     end
 assign n_59 = retime_s3_83_reg_reg_IQ;
 reg retime_s3_84_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_84_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_84_reg_reg_IQ <= n_32;
     end
 assign n_247 = retime_s3_84_reg_reg_IQ;
 reg retime_s3_85_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_85_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_85_reg_reg_IQ <= n_1;
     end
 assign n_17 = retime_s3_85_reg_reg_IQ;
 reg retime_s3_86_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_86_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_86_reg_reg_IQ <= n_82;
     end
 assign n_134 = retime_s3_86_reg_reg_IQ;
 reg retime_s3_88_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_88_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_88_reg_reg_IQ <= n_92;
     end
 assign n_16 = retime_s3_88_reg_reg_IQ;
 reg retime_s3_89_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_89_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_89_reg_reg_IQ <= n_31;
     end
 assign n_15 = retime_s3_89_reg_reg_IQ;
 reg retime_s3_90_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_90_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_90_reg_reg_IQ <= n_140;
     end
 assign n_48 = retime_s3_90_reg_reg_IQ;
 reg retime_s3_91_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_91_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_91_reg_reg_IQ <= n_139;
     end
 assign n_56 = retime_s3_91_reg_reg_IQ;
 reg retime_s3_92_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_92_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_92_reg_reg_IQ <= n_79;
     end
 assign n_116 = retime_s3_92_reg_reg_IQ;
 reg retime_s3_94_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_94_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_94_reg_reg_IQ <= n_0;
     end
 assign n_55 = retime_s3_94_reg_reg_IQ;
 reg retime_s3_99_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_99_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_99_reg_reg_IQ <= n_78;
     end
 assign n_126 = retime_s3_99_reg_reg_IQ;
 reg retime_s3_104_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_104_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_104_reg_reg_IQ <= n_99;
     end
 assign n_52 = retime_s3_104_reg_reg_IQ;
 reg retime_s3_105_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_105_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_105_reg_reg_IQ <= n_30;
     end
 assign n_53 = retime_s3_105_reg_reg_IQ;
 reg retime_s3_106_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_106_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_106_reg_reg_IQ <= n_137;
     end
 assign n_54 = retime_s3_106_reg_reg_IQ;
 reg retime_s3_107_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_107_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_107_reg_reg_IQ <= n_29;
     end
 assign n_127 = retime_s3_107_reg_reg_IQ;
 reg retime_s3_110_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_110_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_110_reg_reg_IQ <= n_77;
     end
 assign n_50 = retime_s3_110_reg_reg_IQ;
 reg retime_s3_111_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_111_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_111_reg_reg_IQ <= n_100;
     end
 assign n_205 = retime_s3_111_reg_reg_IQ;
 reg retime_s3_112_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_112_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_112_reg_reg_IQ <= n_28;
     end
 assign n_60 = retime_s3_112_reg_reg_IQ;
 reg retime_s3_113_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_113_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_113_reg_reg_IQ <= n_27;
     end
 assign n_118 = retime_s3_113_reg_reg_IQ;
 reg retime_s3_114_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_114_reg_reg_IQ <= 1'B1;
     else begin
         retime_s3_114_reg_reg_IQ <= n_26;
     end
 assign n_13 = retime_s3_114_reg_reg_IQ;
 reg retime_s3_116_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_116_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_116_reg_reg_IQ <= n_103;
     end
 assign n_121 = retime_s3_116_reg_reg_IQ;
 reg retime_s3_119_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s3_119_reg_reg_IQ <= 1'B0;
     else begin
         retime_s3_119_reg_reg_IQ <= n_148;
     end
 assign n_128 = retime_s3_119_reg_reg_IQ;
 reg retime_s4_1_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_1_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_1_reg_reg_IQ <= n_75;
     end
 assign n_11 = retime_s4_1_reg_reg_IQ;
 reg retime_s4_2_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_2_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_2_reg_reg_IQ <= n_25;
     end
 assign n_117 = retime_s4_2_reg_reg_IQ;
 reg retime_s4_60_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_60_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_60_reg_reg_IQ <= n_68;
     end
 assign n_9 = retime_s4_60_reg_reg_IQ;
 reg retime_s4_65_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_65_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_65_reg_reg_IQ <= n_34;
     end
 assign n_119 = retime_s4_65_reg_reg_IQ;
 reg retime_s4_76_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_76_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_76_reg_reg_IQ <= n_107;
     end
 assign n_45 = retime_s4_76_reg_reg_IQ;
 reg retime_s4_77_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_77_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_77_reg_reg_IQ <= n_20;
     end
 assign n_44 = retime_s4_77_reg_reg_IQ;
 reg retime_s4_78_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_78_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_78_reg_reg_IQ <= n_189;
     end
 assign n_166 = retime_s4_78_reg_reg_IQ;
 reg retime_s4_79_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_79_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_79_reg_reg_IQ <= n_40;
     end
 assign n_8 = retime_s4_79_reg_reg_IQ;
 reg retime_s4_80_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_80_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_80_reg_reg_IQ <= n_62;
     end
 assign n_113 = retime_s4_80_reg_reg_IQ;
 reg retime_s4_81_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_81_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_81_reg_reg_IQ <= n_112;
     end
 assign n_165 = retime_s4_81_reg_reg_IQ;
 reg retime_s4_82_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_82_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_82_reg_reg_IQ <= n_19;
     end
 assign n_164 = retime_s4_82_reg_reg_IQ;
 reg retime_s4_88_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_88_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_88_reg_reg_IQ <= n_115;
     end
 assign n_161 = retime_s4_88_reg_reg_IQ;
 reg retime_s4_89_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_89_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_89_reg_reg_IQ <= n_18;
     end
 assign n_160 = retime_s4_89_reg_reg_IQ;
 reg retime_s4_90_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_90_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_90_reg_reg_IQ <= n_61;
     end
 assign n_120 = retime_s4_90_reg_reg_IQ;
 reg retime_s4_91_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_91_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_91_reg_reg_IQ <= n_135;
     end
 assign n_7 = retime_s4_91_reg_reg_IQ;
 reg retime_s4_92_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_92_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_92_reg_reg_IQ <= n_125;
     end
 assign n_111 = retime_s4_92_reg_reg_IQ;
 reg retime_s4_93_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_93_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_93_reg_reg_IQ <= n_46;
     end
 assign n_43 = retime_s4_93_reg_reg_IQ;
 reg retime_s4_94_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_94_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_94_reg_reg_IQ <= n_59;
     end
 assign n_42 = retime_s4_94_reg_reg_IQ;
 reg retime_s4_95_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_95_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_95_reg_reg_IQ <= n_247;
     end
 assign n_110 = retime_s4_95_reg_reg_IQ;
 reg retime_s4_96_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_96_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_96_reg_reg_IQ <= n_17;
     end
 assign n_72 = retime_s4_96_reg_reg_IQ;
 reg retime_s4_97_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_97_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_97_reg_reg_IQ <= n_134;
     end
 assign n_41 = retime_s4_97_reg_reg_IQ;
 reg retime_s4_99_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_99_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_99_reg_reg_IQ <= n_16;
     end
 assign n_109 = retime_s4_99_reg_reg_IQ;
 reg retime_s4_100_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_100_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_100_reg_reg_IQ <= n_15;
     end
 assign n_108 = retime_s4_100_reg_reg_IQ;
 reg retime_s4_101_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_101_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_101_reg_reg_IQ <= n_48;
     end
 assign n_6 = retime_s4_101_reg_reg_IQ;
 reg retime_s4_102_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_102_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_102_reg_reg_IQ <= n_56;
     end
 assign n_73 = retime_s4_102_reg_reg_IQ;
 reg retime_s4_109_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_109_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_109_reg_reg_IQ <= n_126;
     end
 assign n_5 = retime_s4_109_reg_reg_IQ;
 reg retime_s4_121_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_121_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_121_reg_reg_IQ <= n_205;
     end
 assign n_106 = retime_s4_121_reg_reg_IQ;
 reg retime_s4_122_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_122_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_122_reg_reg_IQ <= n_60;
     end
 assign n_158 = retime_s4_122_reg_reg_IQ;
 reg retime_s4_123_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_123_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_123_reg_reg_IQ <= n_118;
     end
 assign n_39 = retime_s4_123_reg_reg_IQ;
 reg retime_s4_124_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_124_reg_reg_IQ <= 1'B1;
     else begin
         retime_s4_124_reg_reg_IQ <= n_13;
     end
 assign n_157 = retime_s4_124_reg_reg_IQ;
 reg retime_s4_126_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_126_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_126_reg_reg_IQ <= n_121;
     end
 assign n_122 = retime_s4_126_reg_reg_IQ;
 reg retime_s4_129_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s4_129_reg_reg_IQ <= 1'B0;
     else begin
         retime_s4_129_reg_reg_IQ <= n_128;
     end
 assign n_38 = retime_s4_129_reg_reg_IQ;
 reg retime_s5_1_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_1_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_1_reg_reg_IQ <= n_11;
     end
 assign n_37 = retime_s5_1_reg_reg_IQ;
 reg retime_s5_2_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_2_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_2_reg_reg_IQ <= n_117;
     end
 assign n_4 = retime_s5_2_reg_reg_IQ;
 reg retime_s5_44_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_44_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_44_reg_reg_IQ <= n_44;
     end
 assign n_35 = retime_s5_44_reg_reg_IQ;
 reg retime_s5_45_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_45_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_45_reg_reg_IQ <= n_166;
     end
 assign n_3 = retime_s5_45_reg_reg_IQ;
 reg retime_s5_46_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_46_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_46_reg_reg_IQ <= n_8;
     end
 assign n_98 = retime_s5_46_reg_reg_IQ;
 reg retime_s5_47_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_47_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_47_reg_reg_IQ <= n_113;
     end
 assign n_97 = retime_s5_47_reg_reg_IQ;
 reg retime_s5_55_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_55_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_55_reg_reg_IQ <= n_161;
     end
 assign n_151 = retime_s5_55_reg_reg_IQ;
 reg retime_s5_56_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_56_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_56_reg_reg_IQ <= n_160;
     end
 assign n_95 = retime_s5_56_reg_reg_IQ;
 reg retime_s5_58_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_58_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_58_reg_reg_IQ <= n_7;
     end
 assign n_94 = retime_s5_58_reg_reg_IQ;
 reg retime_s5_59_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_59_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_59_reg_reg_IQ <= n_111;
     end
 assign n_93 = retime_s5_59_reg_reg_IQ;
 reg retime_s5_61_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_61_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_61_reg_reg_IQ <= n_42;
     end
 assign n_2 = retime_s5_61_reg_reg_IQ;
 reg retime_s5_62_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_62_reg_reg_IQ <= 1'B1;
     else begin
         retime_s5_62_reg_reg_IQ <= n_110;
     end
 assign n_91 = retime_s5_62_reg_reg_IQ;
 reg retime_s5_63_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_63_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_63_reg_reg_IQ <= n_72;
     end
 assign n_90 = retime_s5_63_reg_reg_IQ;
 reg retime_s5_66_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_66_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_66_reg_reg_IQ <= n_109;
     end
 assign n_89 = retime_s5_66_reg_reg_IQ;
 reg retime_s5_81_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_81_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_81_reg_reg_IQ <= n_106;
     end
 assign n_147 = retime_s5_81_reg_reg_IQ;
 reg retime_s5_83_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_83_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_83_reg_reg_IQ <= n_39;
     end
 assign n_81 = retime_s5_83_reg_reg_IQ;
 reg retime_s5_86_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_86_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_86_reg_reg_IQ <= n_122;
     end
 assign n_83 = retime_s5_86_reg_reg_IQ;
 reg retime_s5_89_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s5_89_reg_reg_IQ <= 1'B0;
     else begin
         retime_s5_89_reg_reg_IQ <= n_38;
     end
 assign n_143 = retime_s5_89_reg_reg_IQ;
 reg retime_s6_1_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_1_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_1_reg_reg_IQ <= n_37;
     end
 assign n_36 = retime_s6_1_reg_reg_IQ;
 reg retime_s6_2_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_2_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_2_reg_reg_IQ <= n_4;
     end
 assign n_141 = retime_s6_2_reg_reg_IQ;
 reg retime_s6_63_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_63_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_63_reg_reg_IQ <= n_298;
     end
 assign n_145 = retime_s6_63_reg_reg_IQ;
 reg retime_s6_64_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_64_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_64_reg_reg_IQ <= n_296;
     end
 assign n_142 = retime_s6_64_reg_reg_IQ;
 reg retime_s6_66_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_66_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_66_reg_reg_IQ <= n_292;
     end
 assign n_146 = retime_s6_66_reg_reg_IQ;
 reg retime_s6_70_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_70_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_70_reg_reg_IQ <= n_288;
     end
 assign n_149 = retime_s6_70_reg_reg_IQ;
 reg retime_s6_80_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_80_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_80_reg_reg_IQ <= n_3;
     end
 assign n_10 = retime_s6_80_reg_reg_IQ;
 reg retime_s6_82_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_82_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_82_reg_reg_IQ <= n_97;
     end
 assign n_74 = retime_s6_82_reg_reg_IQ;
 reg retime_s6_90_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_90_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_90_reg_reg_IQ <= n_151;
     end
 assign n_71 = retime_s6_90_reg_reg_IQ;
 reg retime_s6_91_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_91_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_91_reg_reg_IQ <= n_95;
     end
 assign n_167 = retime_s6_91_reg_reg_IQ;
 reg retime_s6_92_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_92_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_92_reg_reg_IQ <= n_280;
     end
 assign n_163 = retime_s6_92_reg_reg_IQ;
 reg retime_s6_96_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_96_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_96_reg_reg_IQ <= n_2;
     end
 assign n_69 = retime_s6_96_reg_reg_IQ;
 reg retime_s6_97_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_97_reg_reg_IQ <= 1'B1;
     else begin
         retime_s6_97_reg_reg_IQ <= n_91;
     end
 assign n_173 = retime_s6_97_reg_reg_IQ;
 reg retime_s6_98_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_98_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_98_reg_reg_IQ <= n_90;
     end
 assign n_172 = retime_s6_98_reg_reg_IQ;
 reg retime_s6_99_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_99_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_99_reg_reg_IQ <= n_277;
     end
 assign n_21 = retime_s6_99_reg_reg_IQ;
 reg retime_s6_101_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_101_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_101_reg_reg_IQ <= n_89;
     end
 assign n_175 = retime_s6_101_reg_reg_IQ;
 reg retime_s6_113_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_113_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_113_reg_reg_IQ <= n_147;
     end
 assign n_65 = retime_s6_113_reg_reg_IQ;
 reg retime_s6_114_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_114_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_114_reg_reg_IQ <= n_271;
     end
 assign n_70 = retime_s6_114_reg_reg_IQ;
 reg retime_s6_115_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_115_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_115_reg_reg_IQ <= n_81;
     end
 assign n_177 = retime_s6_115_reg_reg_IQ;
 reg retime_s6_116_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_116_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_116_reg_reg_IQ <= n_269;
     end
 assign n_180 = retime_s6_116_reg_reg_IQ;
 reg retime_s6_118_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_118_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_118_reg_reg_IQ <= n_83;
     end
 assign n_64 = retime_s6_118_reg_reg_IQ;
 reg retime_s6_121_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s6_121_reg_reg_IQ <= 1'B0;
     else begin
         retime_s6_121_reg_reg_IQ <= n_143;
     end
 assign n_104 = retime_s6_121_reg_reg_IQ;
 reg retime_s7_1_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_1_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_1_reg_reg_IQ <= n_36;
     end
 assign n_123 = retime_s7_1_reg_reg_IQ;
 reg retime_s7_2_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_2_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_2_reg_reg_IQ <= n_141;
     end
 assign n_63 = retime_s7_2_reg_reg_IQ;
 reg retime_s7_36_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_36_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_36_reg_reg_IQ <= n_149;
     end
 assign n_132 = retime_s7_36_reg_reg_IQ;
 reg retime_s7_44_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_44_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_44_reg_reg_IQ <= n_10;
     end
 assign n_58 = retime_s7_44_reg_reg_IQ;
 reg retime_s7_52_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_52_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_52_reg_reg_IQ <= n_71;
     end
 assign n_133 = retime_s7_52_reg_reg_IQ;
 reg retime_s7_53_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_53_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_53_reg_reg_IQ <= n_167;
     end
 assign n_57 = retime_s7_53_reg_reg_IQ;
 reg retime_s7_55_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_55_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_55_reg_reg_IQ <= n_69;
     end
 assign n_238 = retime_s7_55_reg_reg_IQ;
 reg retime_s7_56_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_56_reg_reg_IQ <= 1'B1;
     else begin
         retime_s7_56_reg_reg_IQ <= n_173;
     end
 assign n_14 = retime_s7_56_reg_reg_IQ;
 reg retime_s7_57_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_57_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_57_reg_reg_IQ <= n_172;
     end
 assign n_131 = retime_s7_57_reg_reg_IQ;
 reg retime_s7_60_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_60_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_60_reg_reg_IQ <= n_175;
     end
 assign n_129 = retime_s7_60_reg_reg_IQ;
 reg retime_s7_72_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_72_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_72_reg_reg_IQ <= n_65;
     end
 assign n_51 = retime_s7_72_reg_reg_IQ;
 reg retime_s7_77_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s7_77_reg_reg_IQ <= 1'B0;
     else begin
         retime_s7_77_reg_reg_IQ <= n_64;
     end
 assign n_49 = retime_s7_77_reg_reg_IQ;
 reg retime_s8_1_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_1_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_1_reg_reg_IQ <= n_123;
     end
 assign n_47 = retime_s8_1_reg_reg_IQ;
 reg retime_s8_2_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_2_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_2_reg_reg_IQ <= n_63;
     end
 assign n_12 = retime_s8_2_reg_reg_IQ;
 reg retime_s8_85_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_85_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_85_reg_reg_IQ <= n_132;
     end
 assign n_169 = retime_s8_85_reg_reg_IQ;
 reg retime_s8_103_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_103_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_103_reg_reg_IQ <= n_238;
     end
 assign n_170 = retime_s8_103_reg_reg_IQ;
 reg retime_s8_104_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_104_reg_reg_IQ <= 1'B1;
     else begin
         retime_s8_104_reg_reg_IQ <= n_14;
     end
 assign n_168 = retime_s8_104_reg_reg_IQ;
 reg retime_s8_105_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_105_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_105_reg_reg_IQ <= n_131;
     end
 assign n_114 = retime_s8_105_reg_reg_IQ;
 reg retime_s8_108_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s8_108_reg_reg_IQ <= 1'B0;
     else begin
         retime_s8_108_reg_reg_IQ <= n_129;
     end
 assign n_162 = retime_s8_108_reg_reg_IQ;
 reg retime_s9_1_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_1_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_1_reg_reg_IQ <= n_47;
     end
 assign n_176 = retime_s9_1_reg_reg_IQ;
 reg retime_s9_2_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_2_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_2_reg_reg_IQ <= n_12;
     end
 assign n_159 = retime_s9_2_reg_reg_IQ;
 reg retime_s9_36_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_36_reg_reg_IQ <= 1'B0;
     else begin
         retime_s9_36_reg_reg_IQ <= n_290;
     end
 assign n_223 = retime_s9_36_reg_reg_IQ;
 reg retime_s9_54_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s9_54_reg_reg_IQ <= 1'B1;
     else begin
         retime_s9_54_reg_reg_IQ <= n_168;
     end
 assign n_105 = retime_s9_54_reg_reg_IQ;
 assign n_2519 = ~n_2520;
 assign n_2520 = ~n_1456;
 assign n_2521 = ~n_2522;
 assign n_2522 = n_1456;
 assign n_2502 = ~(n_3216 & n_1444);
 assign n_2503 = ~n_1444;
 assign n_2511 = ~n_1449;
 assign n_2516 = ~(n_1456 & {in2[28]});
 assign n_1473 = ~(n_2531 & (~n_1468 | n_1465));
 assign n_2532 = ~n_1465;
 assign n_2536 = ~(n_1470 & n_2532);
 assign n_1502 = (~n_2550 | (n_3237 & n_2553));
 assign n_2542 = ~n_1476;
 assign n_2550 = ~(~n_3192 & n_2554);
 assign n_2531 = ~(n_3229 & n_1465);
 assign n_1500 = ~(n_2551 & (~n_1493 | n_2553));
 assign n_2551 = ~(n_3233 & n_2553);
 assign n_2553 = ~n_2554;
 assign n_2554 = ~n_1489;
 assign n_1513 = ~(n_2565 & (~n_1505 | n_1504));
 assign n_2565 = ~(n_3238 & n_1504);
 assign n_2567 = ~n_1504;
 assign n_1537 = (~n_2581 | (n_3043 & n_1521));
 assign n_1534 = (~n_2580 | (n_3241 & n_1521));
 assign n_1531 = (~n_2583 | (n_1513 & n_1521));
 assign n_1538 = ~((n_2576 | n_2577) & (n_1521 | n_3193));
 assign n_1532 = (~n_2579 | (n_3722 & n_1521));
 assign n_1535 = (~n_2573 | (n_3723 & n_1521));
 assign n_1533 = (~n_2578 | (n_3721 & n_1521));
 assign n_1536 = (~n_2582 | (n_3724 & n_1521));
 assign n_2573 = ~(n_2577 & n_1526);
 assign n_2576 = ~n_3242;
 assign n_2577 = ~n_1521;
 assign n_2578 = ~(n_1524 & n_2577);
 assign n_2579 = ~(n_1523 & n_2577);
 assign n_2580 = ~(n_1525 & n_2577);
 assign n_2581 = ~(n_1528 & n_2577);
 assign n_2582 = ~(n_1527 & n_2577);
 assign n_2583 = ~(n_1522 & n_2577);
 assign n_2590 = ~n_1540;
 assign n_2600 = ~(n_735 & ~n_1540);
 assign n_1579 = ~(n_2602 & (~n_1568 | n_2606));
 assign n_1576 = ~(n_2603 & (~n_1565 | n_2606));
 assign n_1583 = ~(n_2609 & (~n_722 | n_1561));
 assign n_2602 = ~(n_3045 & n_1561);
 assign n_2603 = ~(n_3243 & n_2606);
 assign n_2606 = ~n_2607;
 assign n_2607 = ~n_1561;
 assign n_2609 = ~(n_723 & n_1561);
 assign n_1607 = ~(n_2622 & (~n_1595 | n_1584));
 assign n_2618 = ~(n_3252 & n_2624);
 assign n_2621 = ~(n_3725 & n_2624);
 assign n_2622 = ~(n_1583 & n_1584);
 assign n_2624 = ~n_2623;
 assign n_2623 = ~n_1584;
 assign n_1601 = ~(n_2621 & (~n_1589 | n_2624));
 assign n_1599 = ~(n_2618 & (~n_1587 | n_2624));
 assign n_2637 = ~n_780;
 assign n_1652 = (~n_2652 | (n_2658 & n_1638));
 assign n_2652 = ~(n_3268 & n_2657);
 assign n_2657 = ~n_2658;
 assign n_2658 = ~n_1636;
 assign n_1688 = ~(n_2682 & (~n_1673 | n_1665));
 assign n_1690 = ~(n_2674 & (~n_1675 | n_1665));
 assign n_1692 = ~(n_2673 & (~n_1677 | n_1665));
 assign n_2673 = ~(n_3283 & n_1665);
 assign n_2674 = ~(n_3284 & n_1665);
 assign n_2677 = ~n_1665;
 assign n_2678 = ~(n_618 & n_1665);
 assign n_2682 = ~(n_3277 & n_1665);
 assign n_1695 = ~(n_2678 & (~n_615 | n_1665));
 assign n_2694 = ~(n_1695 & n_1696);
 assign n_2695 = ~(n_3293 & n_1696);
 assign n_2696 = ~n_1696;
 assign n_1725 = ~(n_2695 & (~n_1709 | n_1696));
 assign n_2698 = ~(n_717 & n_1696);
 assign n_1727 = ~(n_2694 & (~n_1711 | n_1696));
 assign n_1728 = ~(n_2698 & (~n_714 | n_1696));
 assign n_2717 = ~n_2719;
 assign n_2719 = ~n_1729;
 assign n_1791 = ~(n_2753 & n_2736);
 assign n_1783 = ~(n_2737 & (~n_1765 | n_2748));
 assign n_1788 = ~(n_2744 & (~n_1770 | n_2748));
 assign n_1799 = ~(n_2738 & (~n_1781 | n_2748));
 assign n_2736 = ~(n_3320 & n_2748);
 assign n_2737 = ~(n_3729 & n_2748);
 assign n_2738 = ~(n_3057 & n_1764);
 assign n_2744 = ~(n_3317 & n_2748);
 assign n_2747 = ~n_1764;
 assign n_2749 = ~n_2748;
 assign n_2748 = n_1764;
 assign n_2753 = ~(n_1773 & n_2747);
 assign n_1828 = ~(n_2775 & (~n_1809 | n_1801));
 assign n_2775 = ~(n_3733 & n_1801);
 assign n_2781 = ~n_1801;
 assign n_2805 = ~n_3699;
 assign n_1916 = ~(n_2826 & (~n_1895 | n_1881));
 assign n_1921 = ~(n_2829 & (~n_1900 | n_1881));
 assign n_2826 = ~(n_3346 & n_1881);
 assign n_2829 = ~(n_3355 & n_1881);
 assign n_2833 = ~n_1881;
 assign n_2863 = ~n_1924;
 assign n_2889 = ~n_1969;
 assign n_2041 = (~n_921 | (n_913 & n_938));
 assign n_2897 = ~(n_300 & n_2017);
 assign n_300 = ~n_2016;
 assign n_2105 = ~(n_2944 & (~n_2080 | n_2065));
 assign n_2108 = ~(n_2947 & (~n_2083 | n_2065));
 assign n_2944 = ~(n_933 & n_2065);
 assign n_2947 = ~(n_931 & n_2065);
 assign n_2949 = ~n_2065;
 assign n_2160 = ~(n_2972 & (~n_2134 | n_2116));
 assign n_2166 = ~(n_2978 & (~n_2140 | n_2116));
 assign n_2972 = ~(n_2108 & n_2116);
 assign n_2978 = ~(n_3060 & n_2116);
 assign n_2979 = ~n_2116;
 assign n_3009 = ~n_2169;
 assign n_2256 = ((n_3493 & n_2224) | (n_3034 & n_2228));
 assign n_2259 = ((n_3494 & n_2224) | (n_3034 & n_2231));
 assign n_2260 = (~n_3030 | (n_3034 & n_2232));
 assign n_2254 = ((n_3504 & n_2224) | (n_3034 & n_2226));
 assign n_2255 = ((n_3505 & n_2224) | (n_3034 & n_2227));
 assign n_2258 = ((n_3507 & n_2224) | (n_3034 & n_2230));
 assign n_3030 = ~(n_3496 & n_2224);
 assign n_3034 = ~n_2224;
 assign n_2328 = ((n_2299 & ~n_3686) | (n_3523 & n_3686));
 assign n_2314 = ((n_2285 & ~n_3686) | (n_2256 & n_3686));
 assign n_2317 = ((n_2288 & ~n_3686) | (n_2259 & n_3686));
 assign n_2324 = ((n_2295 & ~n_3686) | (n_3516 & n_3686));
 assign n_2337 = ((n_2308 & ~n_3686) | (n_3068 & n_3686));
 assign n_2338 = ((n_2309 & ~n_3686) | (n_3517 & n_3686));
 assign n_2339 = ((n_3686 & n_517) | (n_301 & n_515));
 assign n_2318 = ((n_2289 & ~n_3686) | (n_2260 & n_3686));
 assign n_2325 = ((n_2296 & ~n_3686) | (n_3518 & n_3686));
 assign n_2326 = ((n_2297 & ~n_3686) | (n_3519 & n_3686));
 assign n_2315 = ((n_2286 & ~n_3686) | (n_3520 & n_3686));
 assign n_2319 = ((n_2290 & ~n_3686) | (n_3521 & n_3686));
 assign n_2327 = ((n_2298 & ~n_3686) | (n_3522 & n_3686));
 assign n_2311 = ((n_2282 & ~n_3686) | (n_3524 & n_3686));
 assign n_2321 = ((n_3528 & n_3686) | (n_301 & n_2292));
 assign n_2329 = ((n_3535 & n_3686) | (n_301 & n_2300));
 assign n_2312 = ((n_1047 & n_1045) | (n_1024 & n_1046));
 assign n_2313 = ((n_2255 & n_3686) | (n_301 & n_2284));
 assign n_2330 = ((n_3526 & n_3686) | (n_301 & n_2301));
 assign n_2331 = ((n_3527 & n_3686) | (n_301 & n_2302));
 assign n_2316 = ((n_2258 & n_3686) | (n_301 & n_2287));
 assign n_2320 = ((n_3515 & n_3686) | (n_301 & n_2291));
 assign n_2332 = ((n_3529 & n_3686) | (n_301 & n_2303));
 assign n_2322 = ((n_3530 & n_3686) | (n_301 & n_2293));
 assign n_2333 = ((n_3531 & n_3686) | (n_301 & n_2304));
 assign n_2334 = ((n_3532 & n_3686) | (n_301 & n_2305));
 assign n_2323 = ((n_3533 & n_3686) | (n_301 & n_2294));
 assign n_2335 = ((n_3534 & n_3686) | (n_301 & n_2306));
 assign n_2336 = ((n_3525 & n_3686) | (n_301 & n_2307));
 assign n_301 = ~n_3686;
 assign n_2378 = ((n_2348 & ~n_2340) | (n_1019 & n_2340));
 assign n_2374 = ((n_2344 & ~n_2340) | (n_1022 & n_2340));
 assign n_2377 = ((n_2347 & ~n_2340) | (n_1020 & n_2340));
 assign n_2384 = ((n_2354 & ~n_2340) | (n_1017 & n_2340));
 assign n_2397 = ((n_2367 & ~n_2340) | (n_1021 & n_2340));
 assign n_2398 = ((n_2368 & ~n_2340) | (n_1025 & n_2340));
 assign n_2399 = ((n_2369 & ~n_2340) | (n_1026 & n_2340));
 assign n_2371 = ((n_2341 & ~n_2340) | (n_1032 & n_2340));
 assign n_2385 = ((n_2355 & ~n_2340) | (n_1028 & n_2340));
 assign n_2400 = ((n_508 & ~n_2340) | (n_511 & n_2340));
 assign n_2386 = ((n_2356 & ~n_2340) | (n_1029 & n_2340));
 assign n_2375 = ((n_2345 & ~n_2340) | (n_1030 & n_2340));
 assign n_2379 = ((n_2349 & ~n_2340) | (n_1035 & n_2340));
 assign n_2387 = ((n_2357 & ~n_2340) | (n_1031 & n_2340));
 assign n_2388 = ((n_2358 & ~n_2340) | (n_1023 & n_2340));
 assign n_2381 = ((n_2351 & ~n_2340) | (n_1027 & n_2340));
 assign n_2389 = ((n_2359 & ~n_2340) | (n_1036 & n_2340));
 assign n_2372 = ((n_2342 & ~n_2340) | (n_2312 & n_2340));
 assign n_2373 = ((n_2343 & ~n_2340) | (n_1018 & n_2340));
 assign n_2390 = ((n_2360 & ~n_2340) | (n_1034 & n_2340));
 assign n_2391 = ((n_2361 & ~n_2340) | (n_1033 & n_2340));
 assign n_2376 = ((n_2346 & ~n_2340) | (n_1016 & n_2340));
 assign n_2380 = ((n_2350 & ~n_2340) | (n_1037 & n_2340));
 assign n_2392 = ((n_2362 & ~n_2340) | (n_1040 & n_2340));
 assign n_2382 = ((n_2352 & ~n_2340) | (n_1038 & n_2340));
 assign n_2393 = ((n_2363 & ~n_2340) | (n_1039 & n_2340));
 assign n_2394 = ((n_2364 & ~n_2340) | (n_1041 & n_2340));
 assign n_2383 = ((n_2353 & ~n_2340) | (n_1043 & n_2340));
 assign n_2395 = ((n_2365 & ~n_2340) | (n_1042 & n_2340));
 assign n_2396 = ((n_2366 & ~n_2340) | (n_1044 & n_2340));
 assign n_2440 = ((n_2409 & ~n_2401) | (n_1074 & n_2401));
 assign n_2436 = ((n_2405 & ~n_2401) | (n_1087 & n_2401));
 assign n_2439 = ((n_2408 & ~n_2401) | (n_1063 & n_2401));
 assign n_2446 = ((n_2415 & ~n_2401) | (n_1053 & n_2401));
 assign n_2459 = ((n_1076 & ~n_2401) | (n_1071 & n_2401));
 assign n_2460 = ((n_1077 & ~n_2401) | (n_1070 & n_2401));
 assign n_2461 = ((n_1075 & ~n_2401) | (n_1069 & n_2401));
 assign n_2433 = ((n_2402 & ~n_2401) | (n_1068 & n_2401));
 assign n_2447 = ((n_2416 & ~n_2401) | (n_1064 & n_2401));
 assign n_2462 = ((n_1078 & ~n_2401) | (n_1079 & n_2401));
 assign n_2448 = ((n_2417 & ~n_2401) | (n_1060 & n_2401));
 assign n_2463 = ((n_706 & ~n_2401) | (n_1116 & n_2401));
 assign n_2437 = ((n_2406 & ~n_2401) | (n_1105 & n_2401));
 assign n_2441 = ((n_2410 & ~n_2401) | (n_1066 & n_2401));
 assign n_2449 = ((n_1090 & ~n_2401) | (n_1067 & n_2401));
 assign n_2458 = ((n_1100 & ~n_2401) | (n_1102 & n_2401));
 assign n_2442 = ((n_2411 & ~n_2401) | (n_1085 & n_2401));
 assign n_2451 = ((n_1093 & ~n_2401) | (n_1072 & n_2401));
 assign n_2434 = ((n_2403 & ~n_2401) | (n_1073 & n_2401));
 assign n_2435 = ((n_2404 & ~n_2401) | (n_1081 & n_2401));
 assign n_2452 = ((n_1089 & ~n_2401) | (n_1083 & n_2401));
 assign n_2453 = ((n_1095 & ~n_2401) | (n_1080 & n_2401));
 assign n_2438 = ((n_2407 & ~n_2401) | (n_1084 & n_2401));
 assign n_2443 = ((n_2412 & ~n_2401) | (n_1059 & n_2401));
 assign n_2454 = ((n_1094 & ~n_2401) | (n_1048 & n_2401));
 assign n_2444 = ((n_2413 & ~n_2401) | (n_1052 & n_2401));
 assign n_2455 = ((n_1097 & ~n_2401) | (n_1086 & n_2401));
 assign n_2456 = ((n_1098 & ~n_2401) | (n_1088 & n_2401));
 assign n_2445 = ((n_2414 & ~n_2401) | (n_1104 & n_2401));
 assign n_2457 = ((n_1099 & ~n_2401) | (n_1103 & n_2401));
 assign n_2450 = ((n_1092 & ~n_2401) | (n_1058 & n_2401));
 assign in2_95_15_ = ((n_2481 & ~n_2464) | (n_2449 & n_2464));
 assign in2_95_28_ = ((n_2468 & ~n_2464) | (n_2436 & n_2464));
 assign in2_95_25_ = ((n_2471 & ~n_2464) | (n_2439 & n_2464));
 assign in2_95_18_ = ((n_2478 & ~n_2464) | (n_2446 & n_2464));
 assign in2_95_5_ = ((n_2491 & ~n_2464) | (n_2459 & n_2464));
 assign in2_95_4_ = ((n_2492 & ~n_2464) | (n_2460 & n_2464));
 assign in2_95_3_ = ((n_2493 & ~n_2464) | (n_2461 & n_2464));
 assign in2_95_24_ = ((n_2472 & ~n_2464) | (n_2440 & n_2464));
 assign in2_95_17_ = ((n_2479 & ~n_2464) | (n_2447 & n_2464));
 assign in2_95_2_ = ((n_2494 & ~n_2464) | (n_2462 & n_2464));
 assign in2_95_16_ = ((n_2480 & ~n_2464) | (n_2448 & n_2464));
 assign in2_95_1_ = ((n_2495 & ~n_2464) | (n_2463 & n_2464));
 assign in2_95_0_ = ((n_510 & ~n_2464) | (n_1117 & n_2464));
 assign in2_95_27_ = ((n_2469 & ~n_2464) | (n_2437 & n_2464));
 assign in2_95_23_ = ((n_2473 & ~n_2464) | (n_2441 & n_2464));
 assign in2_95_31_ = ((n_2465 & ~n_2464) | (n_2433 & n_2464));
 assign in2_95_6_ = ((n_2490 & ~n_2464) | (n_2458 & n_2464));
 assign in2_95_22_ = ((n_2474 & ~n_2464) | (n_2442 & n_2464));
 assign in2_95_13_ = ((n_2483 & ~n_2464) | (n_2451 & n_2464));
 assign in2_95_30_ = ((n_2466 & ~n_2464) | (n_2434 & n_2464));
 assign in2_95_29_ = ((n_2467 & ~n_2464) | (n_2435 & n_2464));
 assign in2_95_12_ = ((n_2484 & ~n_2464) | (n_2452 & n_2464));
 assign in2_95_11_ = ((n_2485 & ~n_2464) | (n_2453 & n_2464));
 assign in2_95_26_ = ((n_2470 & ~n_2464) | (n_2438 & n_2464));
 assign in2_95_21_ = ((n_2475 & ~n_2464) | (n_2443 & n_2464));
 assign in2_95_10_ = ((n_2486 & ~n_2464) | (n_2454 & n_2464));
 assign in2_95_20_ = ((n_2476 & ~n_2464) | (n_2444 & n_2464));
 assign in2_95_9_ = ((n_2487 & ~n_2464) | (n_2455 & n_2464));
 assign in2_95_8_ = ((n_2488 & ~n_2464) | (n_2456 & n_2464));
 assign in2_95_19_ = ((n_2477 & ~n_2464) | (n_2445 & n_2464));
 assign in2_95_7_ = ((n_2489 & ~n_2464) | (n_2457 & n_2464));
 assign in2_95_14_ = ((n_2482 & ~n_2464) | (n_2450 & n_2464));
 assign n_1441 = ~(n_3720 & (n_3070 & (~n_3689 & ~n_3161)));
 assign n_1444 = ~(sub_181_2_n_29 & sub_181_2_n_30);
 assign sub_181_2_n_30 = ~(sub_181_2_n_28 | (~n_3106 | ~n_3690));
 assign sub_181_2_n_29 = ~(n_3159 | (n_3719 | (n_3689 | n_3161)));
 assign sub_181_2_n_28 = ~((sub_257_2_n_10 & sub_181_2_n_0) | (n_3216 & (sub_257_2_n_10 ^ sub_181_2_n_0)));
 assign n_1445 = ~(sub_181_2_n_0 ^ sub_181_2_n_22);
 assign sub_181_2_n_22 = ({in1[1]} ^ n_3216);
 assign sub_181_2_n_0 = ~(~{in2[30]} & {in1[0]});
 assign sub_200_2_n_5 = ~(~sub_200_2_n_33 | (n_3689 | sub_200_2_n_32));
 assign n_1449 = ~(sub_200_2_n_5 & sub_200_2_n_37);
 assign sub_200_2_n_37 = ~(sub_200_2_n_36 | (~sub_257_2_n_9 | ~n_3537));
 assign sub_200_2_n_36 = ~(sub_200_2_n_0 | (~sub_200_2_n_16 & sub_200_2_n_35));
 assign sub_200_2_n_35 = ~(({in1[1]} & sub_200_2_n_1) | (sub_200_2_n_8 & ({in1[1]} ^ sub_200_2_n_1)));
 assign n_1451 = ~(sub_200_2_n_6 ^ sub_200_2_n_27);
 assign sub_200_2_n_33 = ~(n_3161 | n_3719);
 assign sub_200_2_n_32 = ~(n_3717 & (n_3716 & n_3117));
 assign sub_200_2_n_28 = ~(sub_200_2_n_0 | sub_200_2_n_16);
 assign sub_200_2_n_27 = ({in1[1]} ^ n_3218);
 assign sub_200_2_n_6 = ~sub_200_2_n_1;
 assign sub_200_2_n_16 = ~(~{in1[2]} | n_3217);
 assign sub_200_2_n_8 = ~n_3218;
 assign n_1450 = (sub_200_2_n_35 ^ sub_200_2_n_28);
 assign sub_200_2_n_2 = ~(~{in1[0]} & {in2[29]});
 assign sub_200_2_n_1 = ~({in2[29]} | ~{in1[0]});
 assign sub_200_2_n_0 = ~({in1[2]} | ~n_3217);
 assign n_1456 = ~(sub_219_2_n_44 & (~sub_219_2_n_39 & ~n_3715));
 assign sub_219_2_n_44 = ~(sub_219_2_n_17 & (~sub_219_2_n_3 | n_3538));
 assign n_1457 = ~(sub_219_2_n_29 ^ sub_219_2_n_41);
 assign sub_219_2_n_41 = ~(n_3183 & (sub_219_2_n_38 | sub_219_2_n_9));
 assign sub_219_2_n_39 = ~(n_3720 & sub_219_2_n_26);
 assign sub_219_2_n_37 = ~((sub_257_2_n_10 & sub_219_2_n_4) | (n_3221 & (sub_257_2_n_10 ^ sub_219_2_n_4)));
 assign sub_219_2_n_38 = ~((sub_257_2_n_10 & sub_219_2_n_4) | (n_3221 & (sub_257_2_n_10 ^ sub_219_2_n_4)));
 assign sub_219_2_n_29 = ~(sub_219_2_n_17 & sub_219_2_n_3);
 assign n_1460 = ~(sub_219_2_n_4 & (~{in2[28]} | {in1[0]}));
 assign sub_219_2_n_26 = ~({in1[4]} | ({in1[5]} | ({in1[6]} | {in1[7]})));
 assign sub_219_2_n_17 = ~(~{in1[3]} & n_3219);
 assign sub_219_2_n_9 = ~(~{in1[2]} | n_3220);
 assign n_1458 = (sub_219_2_n_5 ^ sub_219_2_n_38);
 assign sub_219_2_n_5 = ~(n_3183 & ~sub_219_2_n_9);
 assign sub_219_2_n_4 = ~(~{in2[28]} & {in1[0]});
 assign sub_219_2_n_3 = ~({in1[3]} & ~n_3219);
 assign n_1466 = ~(sub_238_2_n_24 ^ sub_238_2_n_36);
 assign n_1465 = ~(sub_238_2_n_38 & sub_238_2_n_28);
 assign sub_238_2_n_38 = ~(n_3164 | (~sub_238_2_n_3 & sub_238_2_n_37));
 assign sub_238_2_n_37 = ~(sub_238_2_n_36 & (~{in1[5]} & ~sub_238_2_n_25));
 assign sub_238_2_n_36 = ~(sub_238_2_n_2 & (~sub_238_2_n_17 | sub_238_2_n_34));
 assign n_1467 = ~(sub_238_2_n_23 ^ sub_238_2_n_33);
 assign sub_238_2_n_34 = ~(sub_238_2_n_16 | (~sub_238_2_n_15 & sub_238_2_n_31));
 assign sub_238_2_n_33 = ~(~sub_238_2_n_16 & (sub_238_2_n_30 | sub_238_2_n_0));
 assign n_1468 = ~((sub_238_2_n_31 & ~sub_238_2_n_4) | (sub_238_2_n_30 & sub_238_2_n_4));
 assign sub_238_2_n_30 = ~sub_238_2_n_31;
 assign sub_238_2_n_31 = ((sub_257_2_n_10 & sub_238_2_n_14) | (n_3224 & (sub_257_2_n_10 ^ sub_238_2_n_14)));
 assign n_1469 = (n_3224 ^ (sub_257_2_n_10 ^ sub_238_2_n_14));
 assign sub_238_2_n_28 = ~({in1[12]} | ({in1[13]} | (~n_3072 | ~sub_238_2_n_26)));
 assign sub_238_2_n_26 = ~({in1[18]} | ({in1[19]} | sub_238_2_n_19));
 assign sub_238_2_n_25 = ~(n_3113 & sub_238_2_n_1);
 assign sub_238_2_n_24 = ~(sub_238_2_n_12 & sub_238_2_n_1);
 assign sub_238_2_n_23 = ~(sub_238_2_n_2 & sub_238_2_n_17);
 assign n_1470 = ~(sub_238_2_n_14 & (~{in2[27]} | {in1[0]}));
 assign sub_238_2_n_19 = ({in1[14]} | ({in1[15]} | ({in1[16]} | {in1[17]})));
 assign sub_238_2_n_17 = ~(sub_238_2_n_9 & {in1[3]});
 assign sub_238_2_n_16 = ~({in1[2]} | sub_238_2_n_8);
 assign sub_238_2_n_15 = ~(~{in1[2]} | n_3229);
 assign sub_238_2_n_14 = ~({in1[0]} & ~{in2[27]});
 assign sub_238_2_n_12 = ~(~{in1[4]} & n_3223);
 assign sub_238_2_n_9 = ~n_3228;
 assign sub_238_2_n_8 = ~n_3229;
 assign sub_257_2_n_10 = ~{in1[1]};
 assign sub_238_2_n_4 = (sub_238_2_n_16 | sub_238_2_n_0);
 assign sub_238_2_n_3 = ~(sub_238_2_n_12 | ({in1[5]} | ~n_3113));
 assign sub_238_2_n_2 = ({in1[3]} | sub_238_2_n_9);
 assign sub_238_2_n_1 = ~(~n_3223 & {in1[4]});
 assign sub_238_2_n_0 = ({in1[2]} & sub_238_2_n_8);
 assign sub_257_2_n_6 = ~({in1[4]} & ~n_3226);
 assign n_1476 = ~(n_708 & (~n_494 & ~n_528));
 assign n_1477 = ~(n_707 ^ n_695);
 assign sub_257_2_n_49 = (~n_3197 | (sub_257_2_n_36 & n_3113));
 assign sub_257_2_n_48 = ~(sub_257_2_n_17 & (~sub_257_2_n_6 | sub_257_2_n_45));
 assign n_1478 = (sub_257_2_n_32 ^ sub_257_2_n_45);
 assign sub_257_2_n_45 = ~sub_257_2_n_44;
 assign sub_257_2_n_44 = ~(sub_257_2_n_2 & (~sub_257_2_n_24 | sub_257_2_n_43));
 assign sub_257_2_n_43 = ~(sub_257_2_n_3 | (~sub_257_2_n_22 & sub_257_2_n_41));
 assign n_1480 = (sub_257_2_n_41 ^ sub_257_2_n_34);
 assign sub_257_2_n_41 = ~(({in1[1]} & sub_257_2_n_16) | (sub_257_2_n_8 & ({in1[1]} ^ sub_257_2_n_16)));
 assign n_1481 = ~(sub_257_2_n_37 ^ sub_257_2_n_25);
 assign sub_257_2_n_39 = ~(n_3072 & (n_3109 & (sub_257_2_n_27 & n_3117)));
 assign sub_257_2_n_37 = ~sub_257_2_n_16;
 assign sub_257_2_n_36 = ~(sub_257_2_n_4 & (sub_257_2_n_17 | sub_257_2_n_18));
 assign sub_257_2_n_35 = ~(sub_257_2_n_6 & sub_257_2_n_19);
 assign sub_257_2_n_34 = ~(sub_257_2_n_3 | sub_257_2_n_1);
 assign sub_257_2_n_33 = ~(sub_257_2_n_4 & sub_257_2_n_19);
 assign sub_257_2_n_32 = ~(sub_257_2_n_17 & sub_257_2_n_6);
 assign sub_257_2_n_31 = ~(sub_257_2_n_2 & sub_257_2_n_24);
 assign n_1482 = ~(sub_257_2_n_37 & (~{in2[26]} | {in1[0]}));
 assign sub_257_2_n_27 = ~({in1[14]} | ({in1[15]} | ({in1[16]} | {in1[17]})));
 assign sub_257_2_n_25 = (~sub_257_2_n_15 | (sub_257_2_n_10 & n_3225));
 assign sub_257_2_n_24 = ~(~sub_257_2_n_9 & sub_257_2_n_11);
 assign sub_257_2_n_22 = ~(~{in1[2]} | n_3231);
 assign sub_257_2_n_19 = ~sub_257_2_n_18;
 assign sub_257_2_n_15 = ~(~sub_257_2_n_10 & sub_257_2_n_8);
 assign sub_257_2_n_18 = ~(~{in1[5]} | n_3230);
 assign sub_257_2_n_17 = ~(~{in1[4]} & n_3226);
 assign sub_257_2_n_16 = ~({in2[26]} | ~{in1[0]});
 assign sub_257_2_n_11 = ~n_1473;
 assign sub_257_2_n_9 = ~{in1[3]};
 assign sub_257_2_n_8 = ~n_3225;
 assign sub_257_2_n_5 = ~(sub_257_2_n_3 | (~sub_257_2_n_1 & sub_257_2_n_41));
 assign sub_257_2_n_4 = ~(~{in1[5]} & n_3230);
 assign sub_257_2_n_3 = ~({in1[2]} | ~n_3231);
 assign sub_257_2_n_2 = ~(sub_257_2_n_9 & ~sub_257_2_n_11);
 assign sub_257_2_n_1 = ~(n_3231 | ~{in1[2]});
 assign n_1479 = (sub_257_2_n_31 ^ sub_257_2_n_5);
 assign sub_276_2_n_4 = ~(sub_276_2_n_26 & ~sub_276_2_n_25);
 assign n_1489 = ~(sub_276_2_n_56 & (~n_3166 & ~n_3165));
 assign n_1490 = ~(sub_276_2_n_4 ^ sub_276_2_n_55);
 assign n_1491 = ~(sub_276_2_n_3 ^ sub_276_2_n_54);
 assign sub_276_2_n_56 = ~(sub_276_2_n_52 & (~sub_276_2_n_36 & ~sub_276_2_n_43));
 assign sub_276_2_n_55 = ~(n_3541 & (~sub_276_2_n_37 | sub_276_2_n_51));
 assign sub_276_2_n_54 = ~(sub_276_2_n_7 & (~sub_276_2_n_24 | sub_276_2_n_51));
 assign n_1492 = (sub_276_2_n_35 ^ sub_276_2_n_51);
 assign sub_276_2_n_52 = ~(~sub_276_2_n_40 & sub_276_2_n_50);
 assign sub_276_2_n_51 = ~sub_276_2_n_50;
 assign sub_276_2_n_50 = ~(sub_276_2_n_1 & (~sub_276_2_n_19 | sub_276_2_n_48));
 assign n_1493 = ~(sub_276_2_n_28 ^ sub_276_2_n_47);
 assign sub_276_2_n_48 = ~(~sub_276_2_n_5 | n_3540);
 assign sub_276_2_n_47 = ~(sub_276_2_n_5 & (sub_276_2_n_6 | sub_276_2_n_17));
 assign n_1494 = (sub_276_2_n_6 ^ sub_276_2_n_2);
 assign sub_276_2_n_43 = ~(~sub_276_2_n_38 | n_3541);
 assign sub_276_2_n_40 = ~(sub_276_2_n_37 & sub_276_2_n_38);
 assign sub_276_2_n_36 = ~(~sub_295_2_n_14 | sub_276_2_n_26);
 assign sub_276_2_n_38 = ~(~sub_295_2_n_14 | sub_276_2_n_25);
 assign sub_276_2_n_37 = ~(sub_276_2_n_23 | sub_276_2_n_18);
 assign sub_276_2_n_35 = ~(sub_276_2_n_7 & sub_276_2_n_24);
 assign n_1496 = ~(sub_276_2_n_16 & (~{in2[25]} | {in1[0]}));
 assign sub_276_2_n_28 = ~(sub_276_2_n_1 & sub_276_2_n_19);
 assign sub_276_2_n_27 = ~(sub_276_2_n_12 ^ n_3237);
 assign sub_276_2_n_24 = ~sub_276_2_n_23;
 assign sub_276_2_n_26 = ~(~n_660 & n_3232);
 assign sub_276_2_n_25 = ~(~n_660 | n_3232);
 assign sub_276_2_n_23 = ~(~n_705 | n_3236);
 assign sub_276_2_n_19 = ~(~sub_276_2_n_9 & sub_276_2_n_11);
 assign sub_276_2_n_18 = ~(~n_642 | n_3235);
 assign sub_276_2_n_17 = ~(~n_425 | n_3234);
 assign sub_276_2_n_16 = ~({in1[0]} & ~{in2[25]});
 assign sub_276_2_n_13 = ~n_425;
 assign sub_276_2_n_12 = ~n_391;
 assign sub_276_2_n_11 = ~n_3233;
 assign sub_276_2_n_9 = ~n_538;
 assign sub_276_2_n_7 = ~(~n_705 & n_3236);
 assign sub_276_2_n_6 = ~((sub_276_2_n_12 & n_644) | (n_3237 & (sub_276_2_n_12 ^ n_644)));
 assign sub_276_2_n_5 = ~(sub_276_2_n_13 & n_3234);
 assign sub_276_2_n_3 = (sub_276_2_n_0 | sub_276_2_n_18);
 assign sub_276_2_n_2 = ~(sub_276_2_n_5 & ~sub_276_2_n_17);
 assign sub_276_2_n_1 = ~(sub_276_2_n_9 & ~sub_276_2_n_11);
 assign sub_276_2_n_0 = ~(n_642 | ~n_3235);
 assign sub_295_2_n_9 = ~(sub_295_2_n_21 & (~sub_295_2_n_49 | sub_295_2_n_3));
 assign n_1505 = (sub_295_2_n_40 ^ sub_295_2_n_62);
 assign n_1504 = ~(sub_295_2_n_59 & (~n_3166 & ~n_3165));
 assign sub_295_2_n_62 = ~(sub_295_2_n_2 | (~sub_295_2_n_30 & sub_295_2_n_58));
 assign n_1506 = ~(sub_295_2_n_7 ^ sub_295_2_n_58);
 assign n_1507 = ~(sub_295_2_n_6 ^ sub_295_2_n_57);
 assign sub_295_2_n_59 = ~(sub_295_2_n_55 & (~sub_295_2_n_32 & ~sub_295_2_n_8));
 assign sub_295_2_n_58 = ~(n_3542 & (~sub_295_2_n_44 | sub_295_2_n_54));
 assign sub_295_2_n_57 = ~(sub_295_2_n_22 & (~sub_295_2_n_29 | sub_295_2_n_54));
 assign n_1508 = (sub_295_2_n_33 ^ sub_295_2_n_54);
 assign sub_295_2_n_55 = ~(~sub_295_2_n_45 & sub_295_2_n_53);
 assign sub_295_2_n_54 = ~sub_295_2_n_53;
 assign sub_295_2_n_53 = ~(sub_295_2_n_0 & (~sub_295_2_n_25 | sub_295_2_n_51));
 assign n_1509 = ~(sub_295_2_n_41 ^ sub_295_2_n_9);
 assign sub_295_2_n_51 = ~(sub_295_2_n_20 | (~sub_295_2_n_16 & sub_295_2_n_49));
 assign n_1510 = ~(sub_295_2_n_49 ^ sub_295_2_n_4);
 assign sub_295_2_n_49 = ((sub_276_2_n_12 & n_487) | (n_3042 & (sub_276_2_n_12 ^ n_487)));
 assign n_1511 = (n_3042 ^ (sub_276_2_n_12 ^ n_487));
 assign sub_295_2_n_45 = ~(sub_295_2_n_44 & sub_295_2_n_39);
 assign sub_295_2_n_43 = ~(sub_295_2_n_2 & sub_295_2_n_24);
 assign sub_295_2_n_41 = ~(sub_295_2_n_0 & sub_295_2_n_25);
 assign sub_295_2_n_40 = ~(sub_295_2_n_31 & sub_295_2_n_24);
 assign sub_295_2_n_44 = ~(sub_295_2_n_28 | sub_295_2_n_10);
 assign n_1512 = ~(sub_295_2_n_19 & (~{in2[24]} | {in1[0]}));
 assign sub_295_2_n_33 = ~(sub_295_2_n_22 & sub_295_2_n_29);
 assign sub_295_2_n_39 = ~(sub_295_2_n_30 | sub_295_2_n_23);
 assign sub_295_2_n_32 = ~sub_295_2_n_31;
 assign sub_295_2_n_29 = ~sub_295_2_n_28;
 assign sub_295_2_n_31 = ~(sub_295_2_n_14 & n_3238);
 assign sub_295_2_n_30 = ~(~n_660 | n_3239);
 assign sub_295_2_n_28 = ~(~n_705 | n_1500);
 assign sub_295_2_n_24 = ~sub_295_2_n_23;
 assign sub_295_2_n_21 = ~sub_295_2_n_20;
 assign sub_295_2_n_25 = ~(sub_295_2_n_13 & n_538);
 assign sub_295_2_n_16 = ~(~n_425 | n_1502);
 assign sub_295_2_n_23 = ~(n_3238 | sub_295_2_n_14);
 assign sub_295_2_n_22 = ~(~n_705 & n_1500);
 assign sub_295_2_n_20 = ~(n_425 | sub_295_2_n_15);
 assign sub_295_2_n_19 = ~({in1[0]} & ~{in2[24]});
 assign sub_295_2_n_15 = ~n_1502;
 assign sub_295_2_n_14 = ~n_683;
 assign sub_295_2_n_13 = ~n_3240;
 assign sub_295_2_n_10 = ~(~n_642 | n_3227);
 assign sub_295_2_n_8 = ~(sub_295_2_n_43 & (~sub_295_2_n_39 | n_3542));
 assign sub_295_2_n_7 = (sub_295_2_n_2 | sub_295_2_n_30);
 assign sub_295_2_n_6 = ~(sub_295_2_n_1 & ~sub_295_2_n_10);
 assign sub_295_2_n_4 = ~(sub_295_2_n_21 & ~sub_295_2_n_3);
 assign sub_295_2_n_3 = (sub_295_2_n_15 & n_425);
 assign sub_295_2_n_2 = ~(n_660 | ~n_3239);
 assign sub_295_2_n_1 = ~(~n_642 & n_3227);
 assign sub_295_2_n_0 = (n_538 | sub_295_2_n_13);
 assign n_1528 = (sub_314_2_n_50 ^ sub_314_2_n_5);
 assign n_1521 = ~(sub_314_2_n_68 & sub_314_2_n_53);
 assign sub_314_2_n_68 = ~(n_3543 & (~sub_314_2_n_45 | sub_314_2_n_67));
 assign sub_314_2_n_67 = ~(sub_314_2_n_64 & (~sub_314_2_n_32 & ~n_401));
 assign n_1522 = (sub_314_2_n_9 ^ sub_314_2_n_10);
 assign n_1523 = (sub_314_2_n_40 ^ sub_314_2_n_63);
 assign sub_314_2_n_64 = ~(~n_3199 & sub_314_2_n_60);
 assign sub_314_2_n_63 = ~(sub_314_2_n_0 | (~sub_314_2_n_22 & sub_314_2_n_58));
 assign n_1524 = ~(sub_314_2_n_7 ^ sub_314_2_n_58);
 assign n_1525 = ~(sub_314_2_n_8 ^ sub_314_2_n_57);
 assign sub_314_2_n_60 = ~(~sub_314_2_n_31 | sub_314_2_n_59);
 assign sub_314_2_n_59 = ~(sub_314_2_n_55 | (~sub_314_2_n_42 | ~sub_314_2_n_41));
 assign sub_314_2_n_58 = ~(sub_314_2_n_44 & (~sub_314_2_n_41 | sub_314_2_n_55));
 assign sub_314_2_n_57 = ~(sub_314_2_n_27 & (~sub_314_2_n_24 | sub_314_2_n_55));
 assign n_1526 = (sub_314_2_n_38 ^ sub_314_2_n_55);
 assign sub_314_2_n_55 = ~(sub_314_2_n_2 | (sub_314_2_n_12 & sub_314_2_n_1));
 assign n_1527 = ~(sub_314_2_n_6 ^ sub_314_2_n_12);
 assign sub_314_2_n_53 = ~(n_614 | (n_456 | sub_314_2_n_52));
 assign sub_314_2_n_52 = ~(sub_314_2_n_48 & (sub_314_2_n_25 & (n_3121 & sub_314_2_n_17)));
 assign sub_314_2_n_50 = ~((sub_276_2_n_12 & n_645) | (n_3242 & (sub_276_2_n_12 ^ n_645)));
 assign sub_314_2_n_48 = ~(~sub_314_2_n_33 | (n_1115 | n_558));
 assign sub_314_2_n_45 = (sub_314_2_n_37 & sub_314_2_n_30);
 assign sub_314_2_n_44 = ~(sub_314_2_n_4 | (n_3200 & sub_314_2_n_29));
 assign sub_314_2_n_40 = ~(sub_314_2_n_31 & sub_314_2_n_21);
 assign sub_314_2_n_42 = ~(sub_314_2_n_22 | sub_314_2_n_20);
 assign sub_314_2_n_41 = ~(sub_314_2_n_23 | sub_314_2_n_28);
 assign sub_314_2_n_39 = ~(sub_276_2_n_12 ^ n_3242);
 assign sub_314_2_n_38 = ~(sub_314_2_n_27 & sub_314_2_n_24);
 assign n_1530 = ~(sub_314_2_n_18 & (~{in2[23]} | {in1[0]}));
 assign sub_314_2_n_35 = ~(sub_314_2_n_0 & sub_314_2_n_21);
 assign sub_314_2_n_33 = ~(n_628 | (n_594 | (n_415 | n_507)));
 assign sub_314_2_n_37 = ~(n_693 | (n_355 | (n_376 | n_527)));
 assign sub_314_2_n_29 = ~sub_314_2_n_28;
 assign sub_314_2_n_27 = ~n_3200;
 assign sub_314_2_n_25 = ~(n_548 | n_670);
 assign sub_314_2_n_32 = ~(~n_445 | n_1513);
 assign sub_314_2_n_31 = ~(~n_683 & n_3722);
 assign sub_314_2_n_30 = ~(n_365 | n_435);
 assign sub_314_2_n_28 = ~(~n_642 | n_3241);
 assign sub_314_2_n_24 = ~sub_314_2_n_23;
 assign sub_314_2_n_21 = ~sub_314_2_n_20;
 assign sub_314_2_n_17 = ~(n_476 | n_568);
 assign sub_314_2_n_23 = ~(~n_705 | n_3723);
 assign sub_314_2_n_22 = ~(~n_660 | n_3721);
 assign sub_314_2_n_20 = ~(~n_683 | n_3722);
 assign sub_314_2_n_19 = ~(~n_425 & n_3043);
 assign sub_314_2_n_18 = ~({in1[0]} & ~{in2[23]});
 assign sub_314_2_n_13 = ~(~n_425 | n_3043);
 assign sub_314_2_n_12 = ~(sub_314_2_n_19 & (sub_314_2_n_50 | sub_314_2_n_13));
 assign sub_314_2_n_10 = ~(sub_314_2_n_59 | (n_3199 | ~sub_314_2_n_31));
 assign sub_314_2_n_9 = (sub_314_2_n_3 | sub_314_2_n_32);
 assign sub_314_2_n_8 = ~(~sub_314_2_n_4 & sub_314_2_n_29);
 assign sub_314_2_n_7 = (sub_314_2_n_0 | sub_314_2_n_22);
 assign sub_314_2_n_6 = ~(~sub_314_2_n_2 & sub_314_2_n_1);
 assign sub_314_2_n_5 = ~(sub_314_2_n_19 & ~sub_314_2_n_13);
 assign sub_314_2_n_4 = ~(n_642 | ~n_3241);
 assign sub_314_2_n_3 = ~(n_445 | ~n_1513);
 assign sub_314_2_n_2 = ~(n_538 | ~n_3724);
 assign sub_314_2_n_1 = ~(~n_3724 & n_538);
 assign sub_314_2_n_0 = ~(n_660 | ~n_3721);
 assign sub_333_2_n_11 = ~(~sub_333_2_n_0 & n_736);
 assign n_1540 = ~(sub_333_2_n_78 & sub_333_2_n_60);
 assign sub_333_2_n_78 = ~(sub_333_2_n_52 & (~sub_333_2_n_43 | sub_333_2_n_76));
 assign n_1541 = (sub_333_2_n_6 ^ sub_333_2_n_75);
 assign sub_333_2_n_76 = ~(n_3169 & (~sub_333_2_n_12 & ~sub_333_2_n_41));
 assign sub_333_2_n_75 = ~(sub_333_2_n_25 | (~sub_333_2_n_12 & n_3169));
 assign n_1542 = ~(sub_333_2_n_10 ^ n_3169);
 assign n_1543 = (sub_333_2_n_11 ^ sub_333_2_n_70);
 assign sub_333_2_n_70 = ~(n_748 | (~n_744 & sub_333_2_n_65));
 assign n_1545 = ~(n_728 ^ sub_333_2_n_67);
 assign n_1544 = ~(sub_333_2_n_9 ^ sub_333_2_n_65);
 assign sub_333_2_n_67 = ~(n_733 & (~n_732 | sub_333_2_n_63));
 assign sub_333_2_n_65 = ~(sub_333_2_n_47 & (~n_739 | sub_333_2_n_63));
 assign n_1546 = (sub_333_2_n_42 ^ sub_333_2_n_63);
 assign sub_333_2_n_63 = ~n_745;
 assign sub_333_2_n_62 = ~(sub_333_2_n_33 & (~n_3194 | sub_333_2_n_58));
 assign n_1547 = ~(n_746 ^ n_730);
 assign sub_333_2_n_60 = ~(n_613 | (n_455 | sub_333_2_n_56));
 assign sub_333_2_n_59 = ~(sub_333_2_n_22 & (sub_333_2_n_55 | sub_333_2_n_4));
 assign sub_333_2_n_58 = ~(sub_333_2_n_21 | (~sub_333_2_n_16 & sub_333_2_n_54));
 assign n_1548 = (n_731 ^ n_729);
 assign sub_333_2_n_56 = ~(sub_333_2_n_49 & (sub_333_2_n_27 & (n_3134 & n_3131)));
 assign sub_333_2_n_55 = ~sub_333_2_n_54;
 assign sub_333_2_n_54 = ((sub_276_2_n_12 & n_576) | (n_3044 & (sub_276_2_n_12 ^ n_576)));
 assign n_1549 = (n_3044 ^ (sub_276_2_n_12 ^ n_576));
 assign sub_333_2_n_52 = ~(sub_333_2_n_48 & (~sub_333_2_n_34 & ~sub_333_2_n_41));
 assign sub_333_2_n_49 = ~(~sub_333_2_n_37 | (n_669 | n_547));
 assign sub_333_2_n_48 = ~(sub_333_2_n_5 & (sub_333_2_n_24 | sub_333_2_n_19));
 assign sub_333_2_n_47 = ~n_741;
 assign sub_333_2_n_46 = ~(sub_333_2_n_2 & (sub_333_2_n_1 | sub_333_2_n_23));
 assign sub_333_2_n_43 = ~(sub_333_2_n_34 | sub_333_2_n_19);
 assign sub_333_2_n_42 = ~(n_733 & n_732);
 assign sub_333_2_n_44 = ~(sub_333_2_n_30 | sub_333_2_n_23);
 assign n_1550 = ~(sub_333_2_n_18 & (~{in2[22]} | {in1[0]}));
 assign sub_333_2_n_37 = ~(n_627 | (n_593 | (n_414 | n_506)));
 assign sub_333_2_n_35 = ~(sub_333_2_n_33 & n_3194);
 assign sub_333_2_n_41 = (n_692 | (n_354 | (n_375 | n_526)));
 assign sub_333_2_n_39 = ~(sub_333_2_n_20 | sub_333_2_n_28);
 assign sub_333_2_n_31 = ~sub_333_2_n_30;
 assign sub_333_2_n_29 = ~sub_333_2_n_28;
 assign sub_333_2_n_27 = ~(n_1114 | n_557);
 assign sub_333_2_n_34 = (n_364 | n_434);
 assign sub_333_2_n_33 = ~(~n_538 & n_1537);
 assign sub_333_2_n_30 = ~(~n_705 | n_1536);
 assign sub_333_2_n_28 = ~(~n_683 | n_1533);
 assign sub_333_2_n_25 = ~sub_333_2_n_24;
 assign sub_333_2_n_22 = ~sub_333_2_n_21;
 assign sub_333_2_n_24 = ~(~n_444 & n_743);
 assign sub_333_2_n_23 = ~(~n_642 | n_1535);
 assign sub_333_2_n_16 = ~(~n_425 | n_1538);
 assign sub_333_2_n_21 = ~(n_425 | sub_333_2_n_14);
 assign sub_333_2_n_20 = ~(~n_660 | n_1534);
 assign sub_333_2_n_19 = ~(~n_400 | n_727);
 assign sub_333_2_n_18 = ~({in1[0]} & ~{in2[22]});
 assign sub_333_2_n_14 = ~n_1538;
 assign sub_333_2_n_12 = ~(~n_444 | n_743);
 assign sub_333_2_n_10 = ~(sub_333_2_n_24 & ~sub_333_2_n_12);
 assign sub_333_2_n_9 = (n_748 | n_744);
 assign sub_333_2_n_8 = ~(sub_333_2_n_2 & ~sub_333_2_n_23);
 assign sub_333_2_n_7 = ~(sub_333_2_n_22 & ~sub_333_2_n_4);
 assign sub_333_2_n_6 = ~(sub_333_2_n_5 & ~sub_333_2_n_19);
 assign sub_333_2_n_5 = ~(~n_400 & n_727);
 assign sub_333_2_n_4 = (n_425 & sub_333_2_n_14);
 assign sub_333_2_n_3 = ~(n_660 | ~n_1534);
 assign sub_333_2_n_2 = ~(~n_642 & n_1535);
 assign sub_333_2_n_1 = ~(~n_705 & n_1536);
 assign sub_333_2_n_0 = ~(n_682 | ~n_738);
 assign n_1570 = (sub_352_2_n_64 ^ sub_352_2_n_10);
 assign n_1561 = ~(n_3172 & sub_352_2_n_86);
 assign n_1562 = (sub_352_2_n_12 ^ sub_352_2_n_16);
 assign n_1563 = (sub_352_2_n_8 ^ sub_352_2_n_84);
 assign sub_352_2_n_86 = (~n_3202 | (sub_352_2_n_65 & n_3129));
 assign n_1565 = (sub_352_2_n_14 ^ sub_352_2_n_81);
 assign sub_352_2_n_84 = ~(sub_352_2_n_28 | (~sub_352_2_n_30 & sub_352_2_n_78));
 assign n_1564 = ~(sub_352_2_n_9 ^ sub_352_2_n_78);
 assign sub_352_2_n_81 = ~(sub_352_2_n_37 | (~sub_352_2_n_43 & sub_352_2_n_15));
 assign n_1566 = ~(sub_352_2_n_54 ^ sub_352_2_n_15);
 assign n_1567 = ~(sub_352_2_n_53 ^ sub_352_2_n_77);
 assign sub_352_2_n_78 = ~(~sub_352_2_n_66 & sub_352_2_n_76);
 assign sub_352_2_n_77 = ~(sub_352_2_n_42 & (~sub_352_2_n_6 | sub_352_2_n_73));
 assign sub_352_2_n_76 = ~(sub_352_2_n_74 & (~sub_352_2_n_51 & ~sub_352_2_n_59));
 assign n_1568 = ~(sub_352_2_n_45 ^ sub_352_2_n_74);
 assign sub_352_2_n_73 = ~sub_352_2_n_74;
 assign sub_352_2_n_74 = ~(sub_352_2_n_2 & (~sub_352_2_n_31 | n_3545));
 assign n_1569 = ~(sub_352_2_n_46 ^ sub_352_2_n_70);
 assign sub_352_2_n_70 = ~(sub_352_2_n_29 & (sub_352_2_n_64 | sub_352_2_n_7));
 assign sub_352_2_n_66 = ~(sub_352_2_n_60 & (sub_352_2_n_13 | sub_352_2_n_51));
 assign sub_352_2_n_65 = ~(sub_352_2_n_57 & (~sub_352_2_n_4 | n_3546));
 assign sub_352_2_n_63 = ~((sub_390_2_n_30 & n_716) | (n_3038 & (sub_390_2_n_30 ^ n_716)));
 assign sub_352_2_n_64 = ~((sub_390_2_n_30 & n_716) | (n_3038 & (sub_390_2_n_30 ^ n_716)));
 assign sub_352_2_n_61 = ~(n_3129 & sub_352_2_n_52);
 assign sub_352_2_n_60 = (~sub_352_2_n_1 & (n_3036 | sub_352_2_n_40));
 assign sub_352_2_n_57 = ~(~n_434 & sub_352_2_n_3);
 assign sub_352_2_n_55 = ~(sub_390_2_n_30 ^ n_3038);
 assign sub_352_2_n_54 = ~(n_3036 & sub_352_2_n_44);
 assign sub_352_2_n_53 = ~(sub_352_2_n_5 & sub_352_2_n_39);
 assign sub_352_2_n_59 = ~(sub_352_2_n_6 & sub_352_2_n_39);
 assign n_1572 = ~(sub_352_2_n_36 & (~{in2[21]} | {in1[0]}));
 assign sub_352_2_n_52 = ~(sub_352_2_n_30 | sub_352_2_n_20);
 assign sub_352_2_n_51 = ~(sub_352_2_n_44 & sub_352_2_n_41);
 assign sub_352_2_n_46 = ~(sub_352_2_n_2 & sub_352_2_n_31);
 assign sub_352_2_n_45 = ~(sub_352_2_n_42 & sub_352_2_n_6);
 assign sub_352_2_n_44 = ~sub_352_2_n_43;
 assign sub_352_2_n_41 = ~sub_352_2_n_40;
 assign sub_352_2_n_39 = ~sub_352_2_n_38;
 assign sub_352_2_n_37 = ~n_3036;
 assign sub_352_2_n_43 = ~(~n_659 | n_3246);
 assign sub_352_2_n_42 = ~(~n_704 & n_3045);
 assign sub_352_2_n_40 = ~(~n_682 | n_3243);
 assign sub_352_2_n_38 = ~(~n_641 | n_3047);
 assign sub_352_2_n_36 = ~({in1[0]} & ~{in2[21]});
 assign sub_352_2_n_28 = ~n_3176;
 assign sub_352_2_n_33 = ~(~n_364 | n_3244);
 assign sub_352_2_n_32 = ~(~n_400 & n_3247);
 assign sub_352_2_n_31 = ~(~sub_352_2_n_23 & sub_352_2_n_22);
 assign sub_352_2_n_27 = ~(~n_424 | n_3248);
 assign sub_352_2_n_30 = ~(~n_444 | n_3249);
 assign sub_352_2_n_29 = ~(~n_424 & n_3248);
 assign sub_352_2_n_23 = ~n_537;
 assign sub_352_2_n_22 = ~n_3245;
 assign sub_352_2_n_20 = ~(~n_400 | n_3247);
 assign n_1571 = ~(n_716 ^ sub_352_2_n_55);
 assign sub_352_2_n_16 = (n_3546 & ~(sub_352_2_n_52 & sub_352_2_n_78));
 assign sub_352_2_n_15 = ~(sub_352_2_n_13 & (sub_352_2_n_59 | sub_352_2_n_73));
 assign sub_352_2_n_14 = ~(~sub_352_2_n_1 & sub_352_2_n_41);
 assign sub_352_2_n_13 = (sub_352_2_n_5 & (sub_352_2_n_42 | sub_352_2_n_38));
 assign sub_352_2_n_12 = (sub_352_2_n_3 | sub_352_2_n_33);
 assign sub_352_2_n_10 = ~(sub_352_2_n_29 & ~sub_352_2_n_7);
 assign sub_352_2_n_9 = ~(n_3176 & ~sub_352_2_n_30);
 assign sub_352_2_n_8 = ~(sub_352_2_n_32 & ~sub_352_2_n_20);
 assign sub_352_2_n_7 = ~(n_3248 | ~n_424);
 assign sub_352_2_n_6 = ~(n_704 & ~n_3045);
 assign sub_352_2_n_5 = ~(~n_641 & n_3047);
 assign sub_352_2_n_4 = ~(n_434 | sub_352_2_n_33);
 assign sub_352_2_n_3 = ~(n_364 | ~n_3244);
 assign sub_352_2_n_2 = ~(sub_352_2_n_23 & ~sub_352_2_n_22);
 assign sub_352_2_n_1 = ~(n_682 | ~n_3243);
 assign n_1595 = ~(n_579 ^ sub_371_2_n_46);
 assign n_1585 = (sub_371_2_n_13 ^ sub_371_2_n_96);
 assign n_1584 = ~(n_3172 & sub_371_2_n_93);
 assign sub_371_2_n_96 = ~(sub_371_2_n_33 | (~sub_371_2_n_36 & sub_371_2_n_14));
 assign n_1587 = (sub_371_2_n_60 ^ sub_371_2_n_92);
 assign n_1586 = ~(sub_371_2_n_11 ^ sub_371_2_n_14);
 assign sub_371_2_n_93 = (~sub_371_2_n_89 | (sub_371_2_n_71 & n_3129));
 assign sub_371_2_n_92 = ~(sub_371_2_n_28 | (~sub_371_2_n_43 & n_3185));
 assign n_1588 = (sub_371_2_n_58 ^ sub_371_2_n_88);
 assign n_1589 = (sub_371_2_n_57 ^ sub_371_2_n_85);
 assign sub_371_2_n_89 = ~(n_3185 & (~sub_371_2_n_52 & ~sub_371_2_n_65));
 assign sub_371_2_n_88 = ~n_3185;
 assign sub_371_2_n_85 = ~(sub_371_2_n_1 | (~sub_371_2_n_40 & sub_371_2_n_15));
 assign n_1590 = ~(sub_371_2_n_12 ^ sub_371_2_n_15);
 assign n_1591 = ~(sub_371_2_n_59 ^ sub_371_2_n_82);
 assign sub_371_2_n_82 = ~(sub_371_2_n_31 & (~sub_371_2_n_6 | sub_371_2_n_79));
 assign sub_371_2_n_81 = ~(sub_371_2_n_78 & (~sub_371_2_n_51 & ~sub_371_2_n_62));
 assign n_1592 = (sub_371_2_n_56 ^ sub_371_2_n_79);
 assign sub_371_2_n_79 = ~sub_371_2_n_78;
 assign sub_371_2_n_78 = ~(sub_371_2_n_8 & (~sub_371_2_n_7 | sub_371_2_n_74));
 assign n_1593 = ~(sub_371_2_n_55 ^ sub_371_2_n_75);
 assign sub_371_2_n_75 = ~(sub_371_2_n_35 & (sub_371_2_n_69 | sub_371_2_n_0));
 assign sub_371_2_n_74 = (~sub_371_2_n_34 & (sub_371_2_n_23 | sub_371_2_n_69));
 assign n_1594 = (sub_371_2_n_69 ^ sub_371_2_n_10);
 assign sub_371_2_n_71 = ~(sub_371_2_n_67 & (~n_3547 & ~sub_371_2_n_4));
 assign sub_371_2_n_70 = (~sub_371_2_n_68 | (sub_371_2_n_1 & sub_371_2_n_39));
 assign sub_371_2_n_69 = ~((sub_390_2_n_30 & n_579) | (n_1583 & (sub_390_2_n_30 ^ n_579)));
 assign sub_371_2_n_68 = ~(sub_371_2_n_64 & sub_371_2_n_61);
 assign sub_371_2_n_67 = ~(sub_371_2_n_63 & n_3548);
 assign sub_371_2_n_65 = ~(n_3129 & n_3548);
 assign sub_371_2_n_64 = ~(sub_371_2_n_5 & (sub_371_2_n_31 | sub_371_2_n_41));
 assign sub_371_2_n_63 = ~(sub_371_2_n_2 & (sub_371_2_n_27 | sub_371_2_n_29));
 assign sub_371_2_n_62 = ~sub_371_2_n_61;
 assign sub_371_2_n_60 = ~(sub_371_2_n_2 & sub_371_2_n_30);
 assign sub_371_2_n_59 = ~(sub_371_2_n_5 & sub_371_2_n_42);
 assign sub_371_2_n_58 = ~(sub_371_2_n_27 & sub_371_2_n_44);
 assign sub_371_2_n_57 = ~(sub_371_2_n_3 & sub_371_2_n_39);
 assign sub_371_2_n_61 = ~(sub_371_2_n_40 | sub_371_2_n_38);
 assign sub_371_2_n_56 = ~(sub_371_2_n_31 & sub_371_2_n_6);
 assign sub_371_2_n_55 = ~(sub_371_2_n_8 & sub_371_2_n_7);
 assign n_1596 = ~(sub_371_2_n_26 & (~{in2[20]} | {in1[0]}));
 assign sub_371_2_n_46 = ~(sub_390_2_n_30 ^ n_1583);
 assign sub_371_2_n_52 = ~(sub_371_2_n_44 & sub_371_2_n_30);
 assign sub_371_2_n_51 = ~(sub_371_2_n_6 & sub_371_2_n_42);
 assign sub_371_2_n_45 = ~sub_371_2_n_3;
 assign sub_371_2_n_44 = ~sub_371_2_n_43;
 assign sub_371_2_n_42 = ~sub_371_2_n_41;
 assign sub_371_2_n_39 = ~sub_371_2_n_38;
 assign sub_371_2_n_43 = ~(~n_444 | n_1576);
 assign sub_371_2_n_41 = ~(~n_641 | n_1579);
 assign sub_371_2_n_40 = ~(~n_659 | n_3253);
 assign sub_371_2_n_38 = ~(~n_682 | n_3725);
 assign sub_371_2_n_35 = ~sub_371_2_n_34;
 assign sub_371_2_n_33 = ~sub_371_2_n_32;
 assign sub_371_2_n_30 = ~sub_371_2_n_29;
 assign sub_371_2_n_28 = ~sub_371_2_n_27;
 assign sub_371_2_n_36 = ~(~n_364 | n_3251);
 assign sub_371_2_n_34 = ~(n_424 | sub_371_2_n_18);
 assign sub_371_2_n_23 = ~(~n_424 | n_3727);
 assign sub_371_2_n_32 = ~(~n_364 & n_3251);
 assign sub_371_2_n_31 = ~(~n_704 & n_3048);
 assign sub_371_2_n_29 = ~(~n_400 | n_3252);
 assign sub_371_2_n_27 = ~(~n_444 & n_1576);
 assign sub_371_2_n_26 = ~({in1[0]} & ~{in2[20]});
 assign sub_371_2_n_21 = ~n_3726;
 assign sub_371_2_n_19 = ~n_364;
 assign sub_371_2_n_18 = ~n_3727;
 assign sub_371_2_n_15 = ~(~sub_371_2_n_64 & (sub_371_2_n_51 | sub_371_2_n_79));
 assign sub_371_2_n_14 = ~(~sub_371_2_n_63 & (sub_371_2_n_52 | sub_371_2_n_88));
 assign sub_371_2_n_13 = (sub_371_2_n_4 | sub_371_2_n_9);
 assign sub_371_2_n_12 = (sub_371_2_n_1 | sub_371_2_n_40);
 assign sub_371_2_n_11 = ~(sub_371_2_n_32 & ~sub_371_2_n_36);
 assign sub_371_2_n_10 = ~(sub_371_2_n_35 & ~sub_371_2_n_0);
 assign sub_371_2_n_9 = ~(n_3250 | ~n_434);
 assign sub_371_2_n_8 = (n_537 | sub_371_2_n_21);
 assign sub_371_2_n_7 = ~(n_537 & sub_371_2_n_21);
 assign sub_371_2_n_6 = ~(n_704 & ~n_3048);
 assign sub_371_2_n_5 = ~(~n_641 & n_1579);
 assign sub_371_2_n_4 = ~(n_434 | ~n_3250);
 assign sub_371_2_n_3 = ~(~n_682 & n_3725);
 assign sub_371_2_n_2 = ~(~n_400 & n_3252);
 assign sub_371_2_n_1 = ~(n_659 | ~n_3253);
 assign sub_371_2_n_0 = (n_424 & sub_371_2_n_18);
 assign sub_390_2_n_21 = (~sub_390_2_n_48 | (sub_390_2_n_46 & sub_390_2_n_17));
 assign n_1611 = ~(n_751 ^ sub_390_2_n_108);
 assign n_1609 = ~(sub_390_2_n_84 & sub_390_2_n_107);
 assign sub_390_2_n_108 = ~(~n_765 & n_771);
 assign sub_390_2_n_107 = ~(sub_390_2_n_11 & (sub_390_2_n_80 & n_3549));
 assign n_1612 = (n_766 ^ n_772);
 assign n_1613 = (n_762 ^ n_769);
 assign n_1610 = ~(n_768 ^ n_764);
 assign sub_390_2_n_103 = ~(~sub_390_2_n_37 & n_3552);
 assign n_1614 = ~(sub_390_2_n_13 ^ sub_390_2_n_96);
 assign n_1615 = (sub_390_2_n_64 ^ sub_390_2_n_21);
 assign sub_390_2_n_98 = ~(~sub_390_2_n_76 & sub_390_2_n_96);
 assign sub_390_2_n_95 = ~(sub_390_2_n_91 & (~sub_390_2_n_0 & ~n_3551));
 assign sub_390_2_n_96 = ~(sub_390_2_n_91 & (~sub_390_2_n_0 & ~n_3551));
 assign n_1616 = ~(sub_390_2_n_57 ^ sub_390_2_n_17);
 assign n_1617 = (sub_390_2_n_65 ^ sub_390_2_n_92);
 assign sub_390_2_n_92 = ~(~sub_390_2_n_55 & sub_390_2_n_88);
 assign sub_390_2_n_91 = ~(sub_390_2_n_87 & (~sub_390_2_n_70 & ~sub_390_2_n_14));
 assign n_1618 = (sub_390_2_n_66 ^ sub_390_2_n_87);
 assign sub_390_2_n_89 = ~(~sub_390_2_n_14 & sub_390_2_n_87);
 assign sub_390_2_n_88 = ~(~sub_390_2_n_35 & sub_390_2_n_87);
 assign sub_390_2_n_87 = ~(sub_390_2_n_85 & sub_390_2_n_4);
 assign n_1619 = ~(sub_390_2_n_56 ^ sub_390_2_n_83);
 assign sub_390_2_n_85 = ~(sub_390_2_n_41 & (~n_3205 | sub_390_2_n_82));
 assign sub_390_2_n_84 = ~(n_1114 | (n_547 | sub_390_2_n_81));
 assign sub_390_2_n_83 = ~(n_3205 & (sub_390_2_n_22 | n_3188));
 assign sub_390_2_n_82 = ~(sub_390_2_n_22 | n_3188);
 assign sub_390_2_n_81 = ~(sub_390_2_n_77 & (sub_390_2_n_44 & (n_3136 & sub_390_2_n_34)));
 assign sub_390_2_n_80 = ~(sub_390_2_n_79 & sub_390_2_n_6);
 assign sub_390_2_n_79 = ~(sub_390_2_n_73 & (~sub_390_2_n_63 | n_3204));
 assign sub_390_2_n_77 = ~(~n_3134 | (n_613 | n_567));
 assign sub_390_2_n_76 = ~(sub_390_2_n_71 & sub_390_2_n_63);
 assign sub_390_2_n_74 = (~sub_390_2_n_3 & (sub_390_2_n_54 | sub_390_2_n_23));
 assign sub_390_2_n_73 = (~sub_390_2_n_5 & (sub_390_2_n_7 | sub_390_2_n_24));
 assign sub_390_2_n_69 = ~(sub_390_2_n_43 | sub_390_2_n_25);
 assign sub_390_2_n_71 = ~(sub_390_2_n_52 | sub_390_2_n_38);
 assign sub_390_2_n_67 = ~(sub_390_2_n_8 | sub_390_2_n_38);
 assign sub_390_2_n_66 = ~(sub_390_2_n_55 | sub_390_2_n_35);
 assign sub_390_2_n_65 = ~(sub_390_2_n_3 | sub_390_2_n_23);
 assign sub_390_2_n_64 = ~(sub_390_2_n_0 | sub_390_2_n_49);
 assign sub_390_2_n_70 = ~(sub_390_2_n_46 & sub_390_2_n_50);
 assign n_1622 = ~(sub_390_2_n_45 & (~{in2[19]} | {in1[0]}));
 assign sub_390_2_n_59 = ~(sub_390_2_n_36 | sub_390_2_n_37);
 assign sub_390_2_n_58 = ~(sub_390_2_n_30 ^ n_3049);
 assign sub_390_2_n_63 = ~(sub_390_2_n_37 | sub_390_2_n_24);
 assign sub_390_2_n_57 = ~(sub_390_2_n_48 & sub_390_2_n_46);
 assign sub_390_2_n_56 = ~(sub_390_2_n_4 & sub_390_2_n_41);
 assign sub_390_2_n_55 = ~sub_390_2_n_54;
 assign sub_390_2_n_53 = ~sub_390_2_n_52;
 assign sub_390_2_n_50 = ~sub_390_2_n_49;
 assign sub_390_2_n_48 = ~sub_390_2_n_47;
 assign sub_390_2_n_44 = ~(n_475 | n_455);
 assign sub_390_2_n_54 = ~(sub_390_2_n_27 & n_3258);
 assign sub_390_2_n_52 = ~(~n_444 | n_1601);
 assign sub_390_2_n_49 = ~(~n_682 | n_3261);
 assign sub_390_2_n_47 = ~(n_659 | sub_390_2_n_28);
 assign sub_390_2_n_46 = ~(sub_390_2_n_28 & n_659);
 assign sub_390_2_n_45 = ~({in1[0]} & ~{in2[19]});
 assign sub_390_2_n_36 = ~sub_390_2_n_7;
 assign sub_390_2_n_35 = ~sub_390_2_n_2;
 assign sub_390_2_n_34 = ~(n_669 | n_557);
 assign sub_390_2_n_43 = (n_375 | n_526);
 assign sub_390_2_n_42 = ~(~n_692 & n_3254);
 assign sub_390_2_n_41 = ~(~sub_352_2_n_23 & sub_390_2_n_31);
 assign sub_390_2_n_38 = ~(~n_400 | n_3255);
 assign sub_390_2_n_37 = ~(~n_364 | n_1599);
 assign sub_390_2_n_31 = ~n_3259;
 assign sub_390_2_n_30 = ~n_390;
 assign sub_390_2_n_28 = ~n_3256;
 assign sub_390_2_n_27 = ~n_704;
 assign sub_390_2_n_25 = ~(~n_692 | n_3254);
 assign sub_390_2_n_24 = ~(~n_434 | n_3260);
 assign sub_390_2_n_23 = ~(~n_641 | n_3257);
 assign sub_390_2_n_22 = ~((sub_390_2_n_30 & n_583) | (n_3049 & (sub_390_2_n_30 ^ n_583)));
 assign n_1620 = (sub_390_2_n_22 ^ sub_390_2_n_9);
 assign sub_390_2_n_19 = ~(sub_390_2_n_98 & ~sub_390_2_n_79);
 assign n_1621 = ~(n_583 ^ sub_390_2_n_58);
 assign sub_390_2_n_17 = ~(sub_390_2_n_74 & sub_390_2_n_89);
 assign sub_390_2_n_14 = ~(sub_390_2_n_2 & ~sub_390_2_n_23);
 assign sub_390_2_n_13 = ~(~sub_390_2_n_1 & sub_390_2_n_53);
 assign sub_390_2_n_12 = (sub_390_2_n_5 | sub_390_2_n_24);
 assign sub_390_2_n_11 = (sub_390_2_n_42 | (sub_390_2_n_43 | n_354));
 assign sub_390_2_n_10 = ~(sub_390_2_n_42 & ~sub_390_2_n_25);
 assign sub_390_2_n_9 = ~(n_3205 & ~n_3188);
 assign sub_390_2_n_8 = ~(n_400 | ~n_3255);
 assign sub_390_2_n_7 = ~(~n_364 & n_1599);
 assign sub_390_2_n_6 = ~(n_354 | (sub_390_2_n_43 | sub_390_2_n_25));
 assign sub_390_2_n_5 = ~(n_434 | ~n_3260);
 assign sub_390_2_n_4 = ~(sub_352_2_n_23 & ~sub_390_2_n_31);
 assign sub_390_2_n_3 = ~(n_641 | ~n_3257);
 assign sub_390_2_n_2 = (sub_390_2_n_27 | n_3258);
 assign sub_390_2_n_1 = ~(n_444 | ~n_1601);
 assign sub_390_2_n_0 = ~(n_682 | ~n_3261);
 assign sub_409_2_n_22 = (~sub_409_2_n_39 | (sub_409_2_n_2 & sub_409_2_n_91));
 assign n_1637 = (sub_409_2_n_16 ^ n_3555);
 assign n_1639 = (sub_409_2_n_65 ^ n_3745);
 assign n_1636 = ~(sub_409_2_n_85 & sub_409_2_n_103);
 assign n_1638 = ~(sub_409_2_n_66 ^ sub_409_2_n_101);
 assign n_1640 = ~(sub_409_2_n_63 ^ n_3554);
 assign n_1641 = ~(sub_409_2_n_17 ^ n_3553);
 assign sub_409_2_n_103 = ~(sub_409_2_n_81 & sub_409_2_n_102);
 assign sub_409_2_n_102 = ~(n_3175 & (~sub_409_2_n_73 & ~sub_409_2_n_72));
 assign sub_409_2_n_101 = ~(~sub_409_2_n_79 & sub_409_2_n_97);
 assign n_1642 = ~(sub_409_2_n_15 ^ n_3175);
 assign n_1643 = ~(sub_409_2_n_10 ^ sub_409_2_n_22);
 assign sub_409_2_n_97 = ~(~sub_409_2_n_73 & n_3175);
 assign n_1644 = ~(sub_409_2_n_54 ^ sub_409_2_n_91);
 assign n_1645 = ~(sub_409_2_n_18 ^ sub_409_2_n_90);
 assign sub_409_2_n_91 = ~(sub_409_2_n_70 & (~sub_409_2_n_60 | sub_409_2_n_88));
 assign sub_409_2_n_90 = ~(sub_409_2_n_24 & (~sub_409_2_n_41 | sub_409_2_n_88));
 assign sub_409_2_n_89 = ~(sub_409_2_n_11 & (~sub_409_2_n_62 & ~sub_409_2_n_61));
 assign sub_409_2_n_88 = ~sub_409_2_n_11;
 assign n_1647 = ~(sub_409_2_n_12 ^ sub_409_2_n_84);
 assign sub_409_2_n_86 = ~(~sub_409_2_n_45 & sub_409_2_n_83);
 assign sub_409_2_n_85 = ~(n_474 | (n_566 | sub_409_2_n_80));
 assign sub_409_2_n_84 = ~(sub_409_2_n_1 & (sub_409_2_n_77 | n_3173));
 assign sub_409_2_n_83 = ~(sub_409_2_n_1 & (sub_409_2_n_77 | n_3173));
 assign n_1648 = (sub_409_2_n_77 ^ sub_409_2_n_9);
 assign sub_409_2_n_81 = ~(sub_409_2_n_75 | (~sub_409_2_n_72 & sub_409_2_n_79));
 assign sub_409_2_n_80 = ~(sub_409_2_n_74 & (sub_409_2_n_46 & (sub_409_2_n_57 & sub_409_2_n_34)));
 assign sub_409_2_n_79 = ~(sub_409_2_n_69 & (~sub_409_2_n_59 | sub_409_2_n_71));
 assign sub_409_2_n_78 = ~(sub_409_2_n_67 & (sub_409_2_n_70 | sub_409_2_n_62));
 assign sub_409_2_n_77 = ~((sub_409_2_n_29 & n_631) | (n_3050 & (sub_409_2_n_29 ^ n_631)));
 assign n_1649 = ~(n_631 ^ sub_409_2_n_55);
 assign sub_409_2_n_75 = ~(sub_409_2_n_42 | (sub_409_2_n_8 & (n_3174 | sub_409_2_n_26)));
 assign sub_409_2_n_74 = ~(~sub_409_2_n_56 | (n_413 | n_592));
 assign sub_409_2_n_73 = ~(sub_409_2_n_68 & sub_409_2_n_59);
 assign sub_409_2_n_72 = ~(sub_409_2_n_53 & (~sub_409_2_n_26 & ~sub_409_2_n_42));
 assign sub_409_2_n_71 = (~sub_409_2_n_4 & (sub_409_2_n_23 | sub_409_2_n_47));
 assign sub_409_2_n_70 = (~sub_409_2_n_7 & (sub_409_2_n_24 | sub_409_2_n_25));
 assign sub_409_2_n_69 = (~sub_409_2_n_5 & (sub_409_2_n_3 | sub_409_2_n_37));
 assign sub_409_2_n_67 = ~(sub_409_2_n_38 & sub_409_2_n_0);
 assign sub_409_2_n_66 = ~(n_3174 & sub_409_2_n_53);
 assign sub_409_2_n_65 = ~(sub_409_2_n_5 | sub_409_2_n_37);
 assign sub_409_2_n_64 = ~(sub_409_2_n_24 & sub_409_2_n_41);
 assign sub_409_2_n_63 = ~(sub_409_2_n_3 & sub_409_2_n_49);
 assign sub_409_2_n_68 = ~(sub_409_2_n_51 | sub_409_2_n_47);
 assign sub_409_2_n_61 = ~sub_409_2_n_60;
 assign n_1650 = ~(sub_409_2_n_35 & (~{in2[18]} | {in1[0]}));
 assign sub_409_2_n_57 = ~(n_484 | (n_602 | (n_342 | n_464)));
 assign sub_409_2_n_56 = ~(n_1113 | (n_546 | (n_668 | n_556)));
 assign sub_409_2_n_62 = ~(sub_409_2_n_2 & sub_409_2_n_0);
 assign sub_409_2_n_60 = ~(sub_409_2_n_40 | sub_409_2_n_25);
 assign sub_409_2_n_59 = ~(sub_409_2_n_48 | sub_409_2_n_37);
 assign sub_409_2_n_55 = ~(sub_409_2_n_29 ^ n_3050);
 assign sub_409_2_n_54 = ~(sub_409_2_n_39 & sub_409_2_n_2);
 assign sub_409_2_n_53 = ~sub_409_2_n_52;
 assign sub_409_2_n_49 = ~sub_409_2_n_48;
 assign sub_409_2_n_46 = ~(n_626 | n_505);
 assign sub_409_2_n_52 = ~(~n_691 | n_3268);
 assign sub_409_2_n_51 = ~(~n_443 | n_3270);
 assign sub_409_2_n_48 = ~(~n_363 | n_3263);
 assign sub_409_2_n_47 = ~(~n_399 | n_3266);
 assign sub_409_2_n_41 = ~sub_409_2_n_40;
 assign sub_409_2_n_39 = ~sub_409_2_n_38;
 assign sub_409_2_n_34 = ~(n_612 | n_454);
 assign sub_409_2_n_45 = ~(~n_536 | n_3271);
 assign sub_409_2_n_44 = ~(~n_536 & n_3271);
 assign sub_409_2_n_43 = ~(n_681 | sub_409_2_n_28);
 assign sub_409_2_n_42 = (n_374 | n_525);
 assign sub_409_2_n_40 = ~(n_3273 | sub_428_2_n_37);
 assign sub_409_2_n_38 = ~(n_658 | sub_409_2_n_31);
 assign sub_409_2_n_37 = ~(~n_433 | n_3269);
 assign sub_409_2_n_35 = ~({in1[0]} & ~{in2[18]});
 assign sub_409_2_n_31 = ~n_3265;
 assign sub_409_2_n_28 = ~n_3264;
 assign sub_409_2_n_26 = ~(~n_353 | n_3262);
 assign sub_409_2_n_25 = ~(~n_640 | n_3267);
 assign sub_409_2_n_24 = ~(sub_428_2_n_37 & n_3273);
 assign sub_409_2_n_23 = ~(sub_428_2_n_41 & n_3270);
 assign n_1646 = (sub_409_2_n_64 ^ sub_409_2_n_88);
 assign sub_409_2_n_18 = (sub_409_2_n_7 | sub_409_2_n_25);
 assign sub_409_2_n_17 = (sub_409_2_n_4 | sub_409_2_n_47);
 assign sub_409_2_n_16 = ~(~sub_409_2_n_8 | sub_409_2_n_26);
 assign sub_409_2_n_15 = ~(sub_409_2_n_23 & ~sub_409_2_n_51);
 assign sub_409_2_n_12 = ~(sub_409_2_n_44 & ~sub_409_2_n_45);
 assign sub_409_2_n_11 = ~(sub_409_2_n_44 & sub_409_2_n_86);
 assign sub_409_2_n_10 = ~(~sub_409_2_n_43 & sub_409_2_n_0);
 assign sub_409_2_n_9 = ~(sub_409_2_n_1 & ~n_3173);
 assign sub_409_2_n_8 = ~(~n_353 & n_3262);
 assign sub_409_2_n_7 = ~(n_640 | ~n_3267);
 assign sub_409_2_n_5 = ~(n_433 | ~n_3269);
 assign sub_409_2_n_4 = ~(n_399 | ~n_3266);
 assign sub_409_2_n_3 = ~(~n_363 & n_3263);
 assign sub_409_2_n_2 = ~(n_658 & sub_409_2_n_31);
 assign sub_409_2_n_1 = ~(~n_423 & n_3272);
 assign sub_409_2_n_0 = ~(n_681 & sub_409_2_n_28);
 assign sub_428_2_n_28 = (~sub_428_2_n_59 | (sub_428_2_n_1 & n_3561));
 assign n_1666 = ~(sub_428_2_n_22 ^ sub_428_2_n_118);
 assign n_1667 = ~(sub_428_2_n_13 ^ sub_428_2_n_117);
 assign n_1669 = ~(sub_428_2_n_19 ^ sub_428_2_n_18);
 assign n_1665 = ~(sub_428_2_n_93 & sub_428_2_n_112);
 assign sub_428_2_n_118 = ~(n_3746 & (~sub_428_2_n_70 | sub_428_2_n_110));
 assign sub_428_2_n_117 = ~(n_3182 & (~sub_428_2_n_50 | sub_428_2_n_110));
 assign n_1668 = ~(sub_428_2_n_71 ^ sub_428_2_n_109);
 assign n_1670 = ~(sub_428_2_n_15 ^ n_3560);
 assign n_1671 = ~(sub_428_2_n_21 ^ n_3556);
 assign sub_428_2_n_113 = ~(~sub_428_2_n_32 & n_3560);
 assign sub_428_2_n_112 = ~(sub_428_2_n_111 & sub_428_2_n_26);
 assign sub_428_2_n_111 = ~(sub_428_2_n_102 & (~sub_428_2_n_81 & ~sub_428_2_n_82));
 assign sub_428_2_n_110 = ~sub_428_2_n_109;
 assign sub_428_2_n_109 = ~(~sub_428_2_n_88 & sub_428_2_n_105);
 assign n_1672 = ~(sub_428_2_n_20 ^ sub_428_2_n_103);
 assign n_1673 = (sub_428_2_n_64 ^ sub_428_2_n_28);
 assign sub_428_2_n_105 = ~(~sub_428_2_n_81 & sub_428_2_n_103);
 assign sub_428_2_n_102 = ~(sub_428_2_n_99 & (~sub_428_2_n_7 & ~n_3558));
 assign sub_428_2_n_103 = ~(sub_428_2_n_99 & (~sub_428_2_n_7 & ~n_3558));
 assign n_1674 = ~(sub_428_2_n_61 ^ n_3561);
 assign n_1675 = (sub_428_2_n_72 ^ n_3562);
 assign sub_428_2_n_99 = ~(sub_428_2_n_95 & (~sub_428_2_n_74 & ~sub_428_2_n_14));
 assign n_1676 = ~(sub_428_2_n_63 ^ sub_428_2_n_95);
 assign sub_428_2_n_95 = ~(sub_428_2_n_0 & (~sub_428_2_n_51 | n_3557));
 assign n_1677 = ~(sub_428_2_n_92 ^ sub_428_2_n_62);
 assign sub_428_2_n_93 = ~(n_342 | (n_464 | sub_428_2_n_89));
 assign sub_428_2_n_92 = ~(sub_428_2_n_4 & (sub_428_2_n_85 | sub_428_2_n_30));
 assign sub_428_2_n_89 = ~(sub_428_2_n_83 & (n_3140 & (n_3139 & n_3138)));
 assign sub_428_2_n_88 = ~(sub_428_2_n_77 & (~sub_428_2_n_76 | sub_428_2_n_80));
 assign sub_428_2_n_87 = ~(sub_428_2_n_12 & (~sub_428_2_n_75 | n_3746));
 assign sub_428_2_n_85 = ~((sub_409_2_n_29 & n_616) | (n_3051 & (sub_409_2_n_29 ^ n_616)));
 assign n_1679 = ~(n_3051 ^ (n_389 ^ n_616));
 assign sub_428_2_n_83 = ~(~n_3141 | (n_1113 | n_556));
 assign sub_428_2_n_82 = ~(sub_428_2_n_70 & sub_428_2_n_75);
 assign sub_428_2_n_81 = ~(n_3559 & sub_428_2_n_76);
 assign sub_428_2_n_80 = (~sub_428_2_n_2 & (sub_428_2_n_57 | sub_428_2_n_34));
 assign sub_428_2_n_78 = (~sub_428_2_n_11 & (sub_428_2_n_43 | sub_428_2_n_31));
 assign sub_428_2_n_77 = (~sub_428_2_n_5 & (n_3180 | sub_428_2_n_33));
 assign sub_428_2_n_72 = ~(sub_428_2_n_11 | sub_428_2_n_31);
 assign sub_428_2_n_76 = ~(sub_428_2_n_32 | sub_428_2_n_33);
 assign sub_428_2_n_75 = ~(sub_428_2_n_52 | n_525);
 assign sub_428_2_n_71 = ~(n_3182 & sub_428_2_n_50);
 assign sub_428_2_n_74 = ~(sub_428_2_n_1 & sub_428_2_n_47);
 assign n_1680 = ~(sub_428_2_n_54 & (~{in2[17]} | {in1[0]}));
 assign sub_428_2_n_64 = ~(sub_428_2_n_7 | sub_428_2_n_46);
 assign sub_428_2_n_63 = ~(sub_428_2_n_8 & sub_428_2_n_29);
 assign sub_428_2_n_62 = ~(sub_428_2_n_0 & sub_428_2_n_51);
 assign sub_428_2_n_70 = ~(sub_428_2_n_49 | sub_428_2_n_48);
 assign sub_428_2_n_61 = ~(sub_428_2_n_59 & sub_428_2_n_1);
 assign sub_428_2_n_59 = ~sub_428_2_n_58;
 assign sub_428_2_n_58 = ~(n_658 | sub_428_2_n_39);
 assign sub_428_2_n_57 = ~(sub_428_2_n_41 & n_3276);
 assign sub_428_2_n_56 = ~(~n_443 | n_3276);
 assign sub_428_2_n_54 = ~({in1[0]} & ~{in2[17]});
 assign sub_428_2_n_50 = ~sub_428_2_n_49;
 assign sub_428_2_n_47 = ~sub_428_2_n_46;
 assign sub_428_2_n_52 = ~(~n_374 | n_3279);
 assign sub_428_2_n_51 = ~(~sub_428_2_n_38 & sub_428_2_n_36);
 assign sub_428_2_n_49 = ~(~n_691 | n_3280);
 assign sub_428_2_n_43 = ~(sub_428_2_n_37 & n_3282);
 assign sub_428_2_n_48 = ~(~n_353 | n_1652);
 assign sub_428_2_n_46 = ~(~n_681 | n_3277);
 assign sub_428_2_n_41 = ~n_443;
 assign sub_428_2_n_40 = ~n_3282;
 assign sub_428_2_n_39 = ~n_3274;
 assign sub_428_2_n_38 = ~n_536;
 assign sub_428_2_n_37 = ~n_703;
 assign sub_428_2_n_36 = ~n_3283;
 assign sub_428_2_n_34 = ~(~n_399 | n_3281);
 assign sub_428_2_n_33 = ~(~n_433 | n_3275);
 assign sub_428_2_n_32 = ~(~n_363 | n_3278);
 assign sub_428_2_n_31 = ~(~n_640 | n_3284);
 assign sub_428_2_n_30 = ~(~n_423 | n_3052);
 assign sub_428_2_n_29 = ~(~sub_428_2_n_37 & sub_428_2_n_40);
 assign n_1678 = (sub_428_2_n_85 ^ sub_428_2_n_17);
 assign sub_428_2_n_26 = ~(sub_428_2_n_87 | (~sub_428_2_n_82 & sub_428_2_n_88));
 assign sub_428_2_n_22 = (sub_428_2_n_6 | sub_428_2_n_52);
 assign sub_428_2_n_21 = (sub_428_2_n_2 | sub_428_2_n_34);
 assign sub_428_2_n_20 = ~(sub_428_2_n_57 & ~sub_428_2_n_56);
 assign sub_428_2_n_19 = (sub_428_2_n_5 | sub_428_2_n_33);
 assign sub_428_2_n_18 = ~(n_3180 & sub_428_2_n_113);
 assign sub_428_2_n_17 = ~(sub_428_2_n_4 & ~sub_428_2_n_30);
 assign sub_428_2_n_15 = ~(n_3180 & ~sub_428_2_n_32);
 assign sub_428_2_n_14 = ~(sub_428_2_n_29 & ~sub_428_2_n_31);
 assign sub_428_2_n_13 = ~(sub_428_2_n_9 & ~sub_428_2_n_48);
 assign sub_428_2_n_12 = ~(sub_428_2_n_6 & ~n_525);
 assign sub_428_2_n_11 = ~(n_640 | ~n_3284);
 assign sub_428_2_n_9 = ~(~n_353 & n_1652);
 assign sub_428_2_n_8 = ~(sub_428_2_n_37 & ~sub_428_2_n_40);
 assign sub_428_2_n_7 = ~(n_681 | ~n_3277);
 assign sub_428_2_n_6 = ~(n_374 | ~n_3279);
 assign sub_428_2_n_5 = ~(n_433 | ~n_3275);
 assign sub_428_2_n_4 = ~(~n_423 & n_3052);
 assign sub_428_2_n_2 = ~(n_399 | ~n_3281);
 assign sub_428_2_n_1 = ~(n_658 & sub_428_2_n_39);
 assign sub_428_2_n_0 = ~(sub_428_2_n_38 & ~sub_428_2_n_36);
 assign sub_447_2_n_23 = (sub_447_2_n_44 | sub_447_2_n_27);
 assign n_1697 = ~(sub_447_2_n_11 ^ sub_447_2_n_139);
 assign sub_447_2_n_139 = ~(sub_447_2_n_50 & (~sub_447_2_n_41 | sub_447_2_n_17));
 assign n_1698 = (sub_447_2_n_82 ^ sub_447_2_n_17);
 assign n_1699 = ~(sub_447_2_n_12 ^ sub_447_2_n_133);
 assign n_1701 = (sub_447_2_n_79 ^ sub_447_2_n_132);
 assign n_1696 = ~sub_447_2_n_134;
 assign sub_447_2_n_134 = ~(sub_447_2_n_107 | (sub_447_2_n_106 & sub_447_2_n_128));
 assign sub_447_2_n_133 = ~(sub_447_2_n_26 & (~sub_447_2_n_43 | n_3189));
 assign sub_447_2_n_132 = ~(sub_447_2_n_1 & (~sub_447_2_n_66 | sub_447_2_n_127));
 assign n_1700 = (sub_447_2_n_80 ^ n_3189);
 assign n_1703 = ~(sub_447_2_n_13 ^ sub_447_2_n_126);
 assign sub_447_2_n_128 = ~(sub_447_2_n_120 & (~sub_447_2_n_92 & ~sub_447_2_n_94));
 assign sub_447_2_n_127 = ~(~sub_447_2_n_91 | sub_447_2_n_123);
 assign sub_447_2_n_126 = ~(sub_447_2_n_6 & (~sub_447_2_n_62 | sub_447_2_n_121));
 assign n_1704 = (sub_447_2_n_69 ^ sub_447_2_n_121);
 assign n_1705 = ~(sub_447_2_n_67 ^ sub_447_2_n_119);
 assign sub_447_2_n_123 = ~(~sub_447_2_n_85 | sub_447_2_n_121);
 assign sub_447_2_n_121 = ~sub_447_2_n_19;
 assign sub_447_2_n_120 = ~(n_3208 & (n_3563 & (sub_447_2_n_111 | sub_447_2_n_23)));
 assign sub_447_2_n_119 = ~(sub_447_2_n_47 & (~sub_447_2_n_58 | sub_447_2_n_116));
 assign n_1706 = ~(sub_447_2_n_68 ^ sub_447_2_n_115);
 assign n_1707 = ~(sub_447_2_n_14 ^ sub_447_2_n_20);
 assign sub_447_2_n_116 = ~(sub_447_2_n_89 | (~sub_447_2_n_23 & n_3713));
 assign sub_447_2_n_115 = ~(~sub_447_2_n_89 & sub_447_2_n_112);
 assign sub_447_2_n_114 = ~(n_3713 & (~sub_447_2_n_76 & ~sub_447_2_n_23));
 assign n_1708 = ~(sub_447_2_n_78 ^ n_3713);
 assign sub_447_2_n_112 = ~(~sub_447_2_n_23 & n_3713);
 assign sub_447_2_n_111 = ~(~sub_447_2_n_76 & sub_447_2_n_109);
 assign sub_447_2_n_109 = ~(sub_447_2_n_25 & (~sub_447_2_n_8 | n_3695));
 assign n_1709 = ~(sub_447_2_n_81 ^ sub_447_2_n_105);
 assign sub_447_2_n_107 = ~(sub_447_2_n_99 & (n_3139 & (n_3138 & sub_447_2_n_55)));
 assign sub_447_2_n_106 = ~(sub_447_2_n_7 | (sub_447_2_n_15 | (sub_447_2_n_16 & sub_447_2_n_93)));
 assign sub_447_2_n_105 = ~(sub_447_2_n_64 & (sub_447_2_n_97 | sub_447_2_n_46));
 assign n_1710 = ~(sub_447_2_n_100 ^ sub_447_2_n_10);
 assign sub_447_2_n_100 = ~sub_447_2_n_97;
 assign sub_447_2_n_99 = ~(n_1113 | (n_556 | (~n_3141 | ~n_3140)));
 assign sub_447_2_n_97 = ~((sub_409_2_n_29 & n_715) | (n_1695 & (sub_409_2_n_29 ^ n_715)));
 assign n_1711 = ~(n_1695 ^ (n_389 ^ n_715));
 assign sub_447_2_n_94 = ~(sub_447_2_n_85 & sub_447_2_n_86);
 assign sub_447_2_n_93 = ~sub_447_2_n_92;
 assign sub_447_2_n_92 = ~(sub_447_2_n_75 & sub_447_2_n_74);
 assign sub_447_2_n_91 = (~sub_447_2_n_2 & (sub_447_2_n_6 | sub_447_2_n_29));
 assign sub_447_2_n_89 = ~sub_447_2_n_88;
 assign sub_447_2_n_88 = (~sub_447_2_n_4 & (sub_447_2_n_24 | sub_447_2_n_27));
 assign sub_447_2_n_87 = (~sub_447_2_n_9 & (sub_447_2_n_1 | sub_447_2_n_30));
 assign sub_447_2_n_84 = ~(sub_447_2_n_0 & sub_447_2_n_49);
 assign sub_447_2_n_86 = ~(sub_447_2_n_65 | sub_447_2_n_30);
 assign sub_447_2_n_82 = ~(sub_447_2_n_50 & sub_447_2_n_41);
 assign sub_447_2_n_81 = ~(sub_447_2_n_25 & n_3207);
 assign sub_447_2_n_80 = ~(sub_447_2_n_26 & sub_447_2_n_43);
 assign sub_447_2_n_79 = ~(sub_447_2_n_9 | sub_447_2_n_30);
 assign sub_447_2_n_78 = ~(sub_447_2_n_24 & sub_447_2_n_45);
 assign sub_447_2_n_85 = ~(sub_447_2_n_61 | sub_447_2_n_29);
 assign sub_447_2_n_77 = ~(sub_447_2_n_1 & sub_447_2_n_66);
 assign n_1712 = ~(sub_447_2_n_56 & (~{in2[16]} | {in1[0]}));
 assign sub_447_2_n_69 = ~(sub_447_2_n_6 & sub_447_2_n_62);
 assign sub_447_2_n_68 = ~(sub_447_2_n_47 & sub_447_2_n_58);
 assign sub_447_2_n_76 = (sub_447_2_n_57 | sub_447_2_n_59);
 assign sub_447_2_n_75 = ~(sub_447_2_n_42 | sub_447_2_n_28);
 assign sub_447_2_n_74 = ~(sub_447_2_n_40 | sub_447_2_n_48);
 assign sub_447_2_n_67 = ~(n_3208 & sub_447_2_n_60);
 assign sub_447_2_n_66 = ~sub_447_2_n_65;
 assign sub_447_2_n_62 = ~sub_447_2_n_61;
 assign sub_447_2_n_60 = ~sub_447_2_n_59;
 assign sub_447_2_n_58 = ~sub_447_2_n_57;
 assign sub_447_2_n_55 = ~(n_342 | n_464);
 assign sub_447_2_n_65 = ~(~n_363 | n_3289);
 assign sub_447_2_n_64 = ~(sub_447_2_n_34 & n_3288);
 assign sub_447_2_n_61 = ~(~n_443 | n_1688);
 assign sub_447_2_n_59 = ~(~n_681 | n_3291);
 assign sub_447_2_n_57 = ~(~n_658 | n_1690);
 assign sub_447_2_n_56 = ~({in1[0]} & ~{in2[16]});
 assign sub_447_2_n_50 = ~sub_447_2_n_0;
 assign sub_447_2_n_49 = ~sub_447_2_n_48;
 assign sub_447_2_n_47 = ~sub_447_2_n_3;
 assign sub_447_2_n_45 = ~sub_447_2_n_44;
 assign sub_447_2_n_43 = ~sub_447_2_n_42;
 assign sub_447_2_n_41 = ~sub_447_2_n_40;
 assign sub_447_2_n_48 = ~(~n_525 | n_3053);
 assign sub_447_2_n_46 = ~(~n_423 | n_3288);
 assign sub_447_2_n_44 = ~(~n_703 | n_1692);
 assign sub_447_2_n_42 = ~(~n_691 | n_3286);
 assign sub_447_2_n_40 = ~(~n_374 | n_3054);
 assign sub_447_2_n_34 = ~n_423;
 assign sub_447_2_n_30 = ~(~n_433 | n_3285);
 assign sub_447_2_n_29 = ~(~n_399 | n_3287);
 assign sub_447_2_n_28 = ~(~n_353 | n_3290);
 assign sub_447_2_n_27 = ~(~n_640 | n_3292);
 assign sub_447_2_n_26 = ~(~n_691 & n_3286);
 assign sub_447_2_n_25 = ~(sub_428_2_n_38 & n_3293);
 assign sub_447_2_n_24 = ~(sub_428_2_n_37 & n_1692);
 assign n_1702 = (sub_447_2_n_77 ^ sub_447_2_n_127);
 assign sub_447_2_n_20 = (~sub_447_2_n_24 | (sub_447_2_n_45 & n_3713));
 assign sub_447_2_n_19 = ~(sub_447_2_n_114 & (n_3208 & n_3563));
 assign sub_447_2_n_17 = ~sub_447_2_n_18;
 assign sub_447_2_n_18 = ~(n_3564 & (~sub_447_2_n_75 | n_3189));
 assign sub_447_2_n_16 = ~(sub_447_2_n_87 & (~sub_447_2_n_86 | sub_447_2_n_91));
 assign sub_447_2_n_15 = ~(sub_447_2_n_84 & (~sub_447_2_n_74 | n_3564));
 assign sub_447_2_n_14 = (sub_447_2_n_4 | sub_447_2_n_27);
 assign sub_447_2_n_13 = (sub_447_2_n_2 | sub_447_2_n_29);
 assign sub_447_2_n_12 = ~(sub_447_2_n_5 & ~sub_447_2_n_28);
 assign sub_447_2_n_11 = ~(~sub_447_2_n_7 & sub_447_2_n_49);
 assign sub_447_2_n_10 = ~(sub_447_2_n_64 & ~sub_447_2_n_46);
 assign sub_447_2_n_9 = ~(n_433 | ~n_3285);
 assign sub_447_2_n_8 = (sub_428_2_n_38 | n_3293);
 assign sub_447_2_n_7 = ~(n_525 | ~n_3053);
 assign sub_447_2_n_6 = ~(~n_443 & n_1688);
 assign sub_447_2_n_5 = ~(~n_353 & n_3290);
 assign sub_447_2_n_4 = ~(n_640 | ~n_3292);
 assign sub_447_2_n_3 = ~(n_658 | ~n_1690);
 assign sub_447_2_n_2 = ~(n_399 | ~n_3287);
 assign sub_447_2_n_1 = ~(~n_363 & n_3289);
 assign sub_447_2_n_0 = ~(n_374 | ~n_3054);
 assign sub_466_2_n_25 = ~(n_703 & ~n_1725);
 assign n_1729 = ~(sub_466_2_n_135 | sub_466_2_n_104);
 assign sub_466_2_n_135 = ~(~sub_466_2_n_93 | sub_466_2_n_129);
 assign n_1732 = (n_3568 ^ sub_466_2_n_66);
 assign n_1733 = (n_829 ^ sub_466_2_n_128);
 assign n_1735 = (n_782 ^ sub_466_2_n_127);
 assign n_1730 = ~(sub_466_2_n_81 ^ sub_466_2_n_123);
 assign sub_466_2_n_129 = ~(sub_466_2_n_123 & (~sub_466_2_n_98 & ~sub_466_2_n_82));
 assign sub_466_2_n_128 = (~n_826 | (sub_466_2_n_122 & n_825));
 assign sub_466_2_n_127 = (~n_819 | (n_3567 & n_816));
 assign n_1734 = ~(sub_466_2_n_77 ^ sub_466_2_n_122);
 assign n_1736 = ~(sub_466_2_n_75 ^ n_3567);
 assign n_1737 = ~(n_814 ^ n_3565);
 assign sub_466_2_n_123 = ~(sub_466_2_n_121 & sub_466_2_n_103);
 assign sub_466_2_n_122 = ~(~sub_466_2_n_97 & sub_466_2_n_117);
 assign sub_466_2_n_121 = ~(n_3171 & (~sub_466_2_n_91 & ~sub_466_2_n_90));
 assign n_1738 = ~(sub_466_2_n_13 ^ n_3171);
 assign n_1739 = (n_803 ^ sub_466_2_n_113);
 assign sub_466_2_n_117 = ~(~sub_466_2_n_90 & n_3171);
 assign sub_466_2_n_113 = (~n_790 | (n_3566 & n_791));
 assign n_1740 = ~(sub_466_2_n_64 ^ n_3566);
 assign n_1741 = (n_823 ^ sub_466_2_n_24);
 assign sub_466_2_n_110 = ~(sub_466_2_n_107 & (~n_824 & ~n_801));
 assign n_1742 = ~(sub_466_2_n_78 ^ sub_466_2_n_107);
 assign sub_466_2_n_107 = ~(n_781 & n_811);
 assign n_1743 = ~(n_810 ^ n_788);
 assign sub_466_2_n_105 = ~(sub_466_2_n_60 & (~sub_466_2_n_53 | sub_466_2_n_100));
 assign sub_466_2_n_104 = ~(sub_466_2_n_5 | (~n_3145 | ~sub_466_2_n_99));
 assign sub_466_2_n_103 = ~(sub_466_2_n_62 | (sub_466_2_n_19 | (sub_466_2_n_97 & sub_466_2_n_92)));
 assign sub_466_2_n_102 = ~(sub_466_2_n_53 & (sub_466_2_n_95 | sub_466_2_n_26));
 assign n_1744 = (sub_466_2_n_16 ^ sub_466_2_n_95);
 assign sub_466_2_n_100 = ~(sub_466_2_n_26 | sub_466_2_n_95);
 assign sub_466_2_n_99 = ~(~n_3144 | (sub_466_2_n_98 | n_565));
 assign sub_466_2_n_98 = ~(n_3143 & (n_3142 & (~n_412 & ~n_591)));
 assign sub_466_2_n_97 = ~(n_818 & (~n_815 | n_817));
 assign sub_466_2_n_96 = ~(n_802 & (n_801 | n_822));
 assign sub_466_2_n_95 = ~((sub_409_2_n_29 & n_491) | (n_1728 & (sub_409_2_n_29 ^ n_491)));
 assign n_1745 = ~(n_1728 ^ (n_389 ^ n_491));
 assign sub_466_2_n_93 = ~(n_565 | ~n_3144);
 assign sub_466_2_n_92 = ~sub_466_2_n_91;
 assign sub_466_2_n_91 = ~(n_798 & n_830);
 assign sub_466_2_n_90 = ~(n_813 & n_815);
 assign sub_466_2_n_89 = (~sub_466_2_n_3 & (sub_466_2_n_9 | sub_466_2_n_50));
 assign sub_466_2_n_88 = (~n_3209 & (sub_466_2_n_1 | n_3190));
 assign sub_466_2_n_87 = ~(~sub_466_2_n_2 | sub_466_2_n_68);
 assign sub_466_2_n_83 = ~(n_797 & n_796);
 assign sub_466_2_n_82 = ~(n_3145 & sub_466_2_n_61);
 assign sub_466_2_n_81 = ~(sub_466_2_n_5 & sub_466_2_n_61);
 assign sub_466_2_n_80 = ~(sub_466_2_n_4 & n_796);
 assign sub_466_2_n_79 = ~(sub_466_2_n_7 | sub_466_2_n_47);
 assign sub_466_2_n_86 = ~(sub_466_2_n_0 & sub_466_2_n_48);
 assign sub_466_2_n_78 = ~(n_808 & n_807);
 assign sub_466_2_n_85 = ~(sub_466_2_n_45 | sub_466_2_n_50);
 assign sub_466_2_n_77 = ~(n_826 & n_825);
 assign sub_466_2_n_76 = ~(sub_466_2_n_3 | sub_466_2_n_50);
 assign sub_466_2_n_75 = ~(n_819 & n_816);
 assign sub_466_2_n_74 = ~(n_3209 | n_3190);
 assign sub_466_2_n_84 = ~(sub_466_2_n_57 | sub_466_2_n_56);
 assign n_1746 = ~(sub_466_2_n_52 & (~{in2[15]} | {in1[0]}));
 assign sub_466_2_n_68 = ~(sub_466_2_n_39 | sub_466_2_n_56);
 assign sub_466_2_n_67 = ~(sub_466_2_n_54 & sub_466_2_n_48);
 assign sub_466_2_n_73 = ~(sub_466_2_n_49 | sub_466_2_n_43);
 assign sub_466_2_n_66 = ~(n_797 | n_784);
 assign sub_466_2_n_65 = ~(sub_466_2_n_10 & sub_466_2_n_60);
 assign sub_466_2_n_64 = ~(n_790 & n_791);
 assign sub_466_2_n_71 = ~(sub_466_2_n_41 | sub_466_2_n_40);
 assign sub_466_2_n_62 = ~sub_466_2_n_4;
 assign sub_466_2_n_58 = ~sub_466_2_n_57;
 assign sub_466_2_n_55 = ~sub_466_2_n_54;
 assign sub_466_2_n_63 = ~(sub_466_2_n_29 & n_3294);
 assign sub_466_2_n_61 = ~(sub_466_2_n_31 & n_473);
 assign sub_466_2_n_60 = ~(~sub_428_2_n_38 & sub_466_2_n_35);
 assign sub_466_2_n_57 = ~(~n_691 | n_3299);
 assign sub_466_2_n_56 = ~(~n_353 | n_3295);
 assign sub_466_2_n_54 = ~(n_658 | sub_466_2_n_34);
 assign sub_466_2_n_53 = ~(sub_447_2_n_34 & n_1727);
 assign sub_466_2_n_52 = ~({in1[0]} & ~{in2[15]});
 assign sub_466_2_n_48 = ~sub_466_2_n_47;
 assign sub_466_2_n_46 = ~sub_466_2_n_45;
 assign sub_466_2_n_44 = ~sub_466_2_n_43;
 assign sub_466_2_n_50 = ~(~n_433 | n_3300);
 assign sub_466_2_n_49 = ~(~n_374 | n_3303);
 assign sub_466_2_n_47 = ~(~n_681 | n_3301);
 assign sub_466_2_n_45 = ~(~n_363 | n_3296);
 assign sub_466_2_n_43 = ~(~n_525 | n_3302);
 assign sub_466_2_n_41 = ~(~n_443 | n_3304);
 assign sub_466_2_n_40 = ~(~n_399 | n_3294);
 assign sub_466_2_n_36 = ~(n_3294 | sub_466_2_n_29);
 assign sub_466_2_n_39 = ~(~n_691 & n_3299);
 assign sub_466_2_n_35 = ~n_3297;
 assign sub_466_2_n_34 = ~n_3305;
 assign sub_409_2_n_29 = ~n_389;
 assign sub_466_2_n_31 = ~n_806;
 assign sub_466_2_n_29 = ~n_399;
 assign sub_466_2_n_26 = ~(~n_423 | n_1727);
 assign sub_466_2_n_24 = (~n_808 | (n_807 & sub_466_2_n_107));
 assign sub_466_2_n_19 = ~(sub_466_2_n_83 & (~n_798 | n_831));
 assign sub_466_2_n_17 = (sub_466_2_n_63 & (sub_466_2_n_8 | sub_466_2_n_36));
 assign sub_466_2_n_16 = ~(sub_466_2_n_53 & ~sub_466_2_n_26);
 assign sub_466_2_n_15 = ~(~sub_466_2_n_2 | sub_466_2_n_56);
 assign sub_466_2_n_14 = ~(sub_466_2_n_25 & ~n_3190);
 assign sub_466_2_n_13 = ~(n_793 & ~n_792);
 assign sub_466_2_n_12 = ~(sub_466_2_n_63 & ~sub_466_2_n_40);
 assign sub_466_2_n_10 = ~(sub_428_2_n_38 & ~sub_466_2_n_35);
 assign sub_466_2_n_9 = ~(~n_363 & n_3296);
 assign sub_466_2_n_8 = ~(~n_443 & n_3304);
 assign sub_466_2_n_7 = ~(n_681 | ~n_3301);
 assign sub_466_2_n_6 = ~(n_374 | ~n_3303);
 assign sub_466_2_n_5 = (n_473 | sub_466_2_n_31);
 assign sub_466_2_n_4 = ~(~n_524 & n_800);
 assign sub_466_2_n_3 = ~(n_433 | ~n_3300);
 assign sub_466_2_n_2 = ~(~n_353 & n_3295);
 assign sub_466_2_n_1 = ~(~n_703 & n_1725);
 assign sub_466_2_n_0 = ~(n_658 & sub_466_2_n_34);
 assign n_1766 = (sub_485_2_n_13 ^ sub_485_2_n_122);
 assign n_1767 = (sub_485_2_n_15 ^ sub_485_2_n_133);
 assign n_1764 = ~(n_3571 | (sub_485_2_n_21 & sub_485_2_n_128));
 assign n_1765 = ~(sub_485_2_n_16 ^ sub_485_2_n_129);
 assign sub_485_2_n_133 = ~(sub_485_2_n_39 | (sub_485_2_n_22 & sub_485_2_n_1));
 assign n_1768 = ~(sub_485_2_n_14 ^ sub_485_2_n_22);
 assign n_1769 = ~(sub_485_2_n_62 ^ sub_485_2_n_127);
 assign n_1771 = (sub_485_2_n_19 ^ sub_485_2_n_126);
 assign sub_485_2_n_129 = ~(sub_485_2_n_56 & (sub_485_2_n_122 | sub_485_2_n_11));
 assign sub_485_2_n_128 = ~(sub_485_2_n_122 | (~sub_485_2_n_93 | ~sub_485_2_n_77));
 assign sub_485_2_n_127 = ~(sub_485_2_n_49 & (~n_3211 | sub_485_2_n_24));
 assign sub_485_2_n_126 = ~(sub_485_2_n_34 | (~sub_485_2_n_33 & sub_485_2_n_121));
 assign n_1770 = (sub_485_2_n_74 ^ sub_485_2_n_24);
 assign n_1772 = (sub_485_2_n_121 ^ sub_485_2_n_63);
 assign n_1773 = ~(sub_485_2_n_20 ^ sub_485_2_n_120);
 assign sub_485_2_n_122 = ~(sub_485_2_n_103 | (~sub_485_2_n_87 & sub_485_2_n_117));
 assign sub_485_2_n_121 = ~(sub_485_2_n_84 & (~sub_485_2_n_72 | sub_485_2_n_116));
 assign sub_485_2_n_120 = ~(sub_485_2_n_45 & (~sub_485_2_n_41 | sub_485_2_n_116));
 assign n_1774 = (sub_485_2_n_60 ^ sub_485_2_n_116);
 assign n_1775 = ~(sub_485_2_n_18 ^ n_3569);
 assign sub_485_2_n_117 = ~(~sub_485_2_n_88 | sub_485_2_n_115);
 assign sub_485_2_n_115 = ~(sub_485_2_n_108 | (~sub_485_2_n_6 | ~n_3572));
 assign sub_485_2_n_116 = ~(sub_485_2_n_108 | (~sub_485_2_n_6 | ~n_3572));
 assign n_1776 = ~(sub_485_2_n_73 ^ sub_485_2_n_110);
 assign n_1777 = ~(sub_485_2_n_17 ^ n_3570);
 assign sub_485_2_n_110 = ~(sub_485_2_n_83 & (~sub_485_2_n_71 | n_3210));
 assign sub_485_2_n_108 = ~(n_3210 | (~sub_485_2_n_79 | ~sub_485_2_n_71));
 assign n_1778 = (sub_485_2_n_76 ^ n_3210);
 assign n_1779 = ~(sub_485_2_n_61 ^ sub_485_2_n_102);
 assign sub_485_2_n_104 = ~(~sub_485_2_n_4 & sub_485_2_n_100);
 assign sub_485_2_n_103 = ~(sub_485_2_n_94 & (~sub_485_2_n_43 & ~sub_485_2_n_91));
 assign sub_485_2_n_102 = ~(~sub_485_2_n_4 & (sub_485_2_n_98 | sub_485_2_n_35));
 assign n_1780 = (sub_485_2_n_97 ^ sub_485_2_n_75);
 assign sub_485_2_n_100 = ~(~sub_485_2_n_35 & sub_485_2_n_97);
 assign sub_485_2_n_98 = ~sub_485_2_n_97;
 assign sub_485_2_n_97 = ((sub_485_2_n_27 & n_404) | (n_3057 & (sub_485_2_n_27 ^ n_404)));
 assign n_1781 = (n_3057 ^ (sub_485_2_n_27 ^ n_404));
 assign sub_485_2_n_95 = ~(sub_485_2_n_93 & n_3145);
 assign sub_485_2_n_94 = ~(sub_485_2_n_92 & sub_485_2_n_88);
 assign sub_485_2_n_93 = ~(n_412 | (n_591 | (~n_3143 | ~n_3142)));
 assign sub_485_2_n_92 = ~(sub_485_2_n_86 & (~sub_485_2_n_78 | sub_485_2_n_84));
 assign sub_485_2_n_91 = ~(sub_485_2_n_66 & (n_3573 | sub_485_2_n_70));
 assign sub_485_2_n_88 = ~(sub_485_2_n_80 | sub_485_2_n_70);
 assign sub_485_2_n_87 = ~(sub_485_2_n_72 & sub_485_2_n_78);
 assign sub_485_2_n_86 = (~sub_485_2_n_5 & (sub_485_2_n_3 | sub_485_2_n_46));
 assign sub_485_2_n_85 = ~(sub_485_2_n_7 & (sub_485_2_n_56 | sub_485_2_n_50));
 assign sub_485_2_n_84 = (~sub_485_2_n_12 & (sub_485_2_n_45 | sub_485_2_n_38));
 assign sub_485_2_n_83 = ~sub_485_2_n_82;
 assign sub_485_2_n_82 = ~(sub_485_2_n_10 & (sub_485_2_n_8 | sub_485_2_n_54));
 assign sub_485_2_n_77 = ~(~n_3145 | sub_485_2_n_11);
 assign sub_485_2_n_80 = ~(n_3211 & sub_485_2_n_52);
 assign sub_485_2_n_79 = ~(sub_485_2_n_47 | sub_485_2_n_55);
 assign sub_485_2_n_76 = ~(sub_485_2_n_8 & sub_485_2_n_37);
 assign sub_485_2_n_75 = ~(sub_485_2_n_4 | sub_485_2_n_35);
 assign sub_485_2_n_78 = ~(sub_485_2_n_33 | sub_485_2_n_46);
 assign sub_485_2_n_74 = ~(sub_485_2_n_49 & n_3211);
 assign sub_485_2_n_73 = ~(sub_485_2_n_0 & sub_485_2_n_48);
 assign sub_485_2_n_66 = ~(sub_485_2_n_39 & sub_485_2_n_42);
 assign n_1782 = ~(sub_485_2_n_32 & (~{in2[14]} | {in1[0]}));
 assign sub_485_2_n_63 = ~(sub_485_2_n_34 | sub_485_2_n_33);
 assign sub_485_2_n_62 = ~(sub_485_2_n_2 & sub_485_2_n_52);
 assign sub_485_2_n_72 = ~(sub_485_2_n_40 | sub_485_2_n_38);
 assign sub_485_2_n_61 = ~(sub_485_2_n_58 & sub_485_2_n_9);
 assign sub_485_2_n_71 = ~(sub_485_2_n_36 | sub_485_2_n_54);
 assign sub_485_2_n_70 = ~(sub_485_2_n_1 & sub_485_2_n_42);
 assign sub_485_2_n_60 = ~(sub_485_2_n_45 & sub_485_2_n_41);
 assign sub_485_2_n_52 = ~sub_485_2_n_51;
 assign sub_485_2_n_48 = ~sub_485_2_n_47;
 assign sub_485_2_n_58 = ~(sub_485_2_n_31 & n_3055);
 assign sub_485_2_n_56 = ~(~n_473 & n_3731);
 assign sub_485_2_n_55 = ~(~n_680 | n_3318);
 assign sub_485_2_n_54 = ~(~n_639 | n_3730);
 assign sub_485_2_n_51 = ~(~n_352 | n_3312);
 assign sub_485_2_n_50 = ~(~n_565 | n_3729);
 assign sub_485_2_n_49 = ~(~n_690 & n_3317);
 assign sub_485_2_n_47 = ~(~n_657 | n_3319);
 assign sub_485_2_n_46 = ~(~n_432 | n_3309);
 assign sub_485_2_n_45 = ~(~n_442 & n_3314);
 assign sub_485_2_n_41 = ~sub_485_2_n_40;
 assign sub_485_2_n_37 = ~sub_485_2_n_36;
 assign sub_485_2_n_34 = ~sub_485_2_n_3;
 assign sub_485_2_n_43 = ~(n_524 | sub_485_2_n_30);
 assign sub_485_2_n_42 = ~(sub_485_2_n_30 & n_524);
 assign sub_485_2_n_40 = ~(~n_442 | n_3314);
 assign sub_485_2_n_39 = ~(n_373 | sub_485_2_n_28);
 assign sub_485_2_n_38 = ~(~n_398 | n_3320);
 assign sub_485_2_n_36 = ~(~n_702 | n_3728);
 assign sub_485_2_n_35 = ~(~n_422 | n_3056);
 assign sub_485_2_n_33 = ~(~n_362 | n_3307);
 assign sub_485_2_n_32 = ~({in1[0]} & ~{in2[14]});
 assign sub_485_2_n_31 = ~n_535;
 assign sub_485_2_n_30 = ~n_3316;
 assign sub_485_2_n_28 = ~n_3308;
 assign sub_485_2_n_27 = ~n_388;
 assign sub_485_2_n_24 = (~sub_485_2_n_92 & (sub_485_2_n_87 | sub_485_2_n_116));
 assign sub_485_2_n_22 = ~(n_3573 & (sub_485_2_n_80 | sub_485_2_n_24));
 assign sub_485_2_n_21 = ~(~n_3144 | sub_485_2_n_50);
 assign sub_485_2_n_20 = (sub_485_2_n_12 | sub_485_2_n_38);
 assign sub_485_2_n_19 = (sub_485_2_n_5 | sub_485_2_n_46);
 assign sub_485_2_n_18 = ~(sub_485_2_n_6 & ~sub_485_2_n_55);
 assign sub_485_2_n_17 = ~(sub_485_2_n_10 & ~sub_485_2_n_54);
 assign sub_485_2_n_16 = ~(sub_485_2_n_7 & ~sub_485_2_n_50);
 assign sub_485_2_n_15 = ~(~sub_485_2_n_43 & sub_485_2_n_42);
 assign sub_485_2_n_14 = ~(~sub_485_2_n_39 & sub_485_2_n_1);
 assign sub_485_2_n_13 = ~(sub_485_2_n_56 & ~sub_485_2_n_11);
 assign sub_485_2_n_12 = ~(n_398 | ~n_3320);
 assign sub_485_2_n_11 = ~(n_3731 | ~n_473);
 assign sub_485_2_n_10 = ~(~n_639 & n_3730);
 assign sub_485_2_n_9 = (sub_485_2_n_31 | n_3055);
 assign sub_485_2_n_8 = ~(~n_702 & n_3728);
 assign sub_485_2_n_7 = ~(~n_565 & n_3729);
 assign sub_485_2_n_6 = ~(~n_680 & n_3318);
 assign sub_485_2_n_5 = ~(n_432 | ~n_3309);
 assign sub_485_2_n_4 = ~(n_422 | ~n_3056);
 assign sub_485_2_n_3 = ~(~n_362 & n_3307);
 assign sub_485_2_n_2 = ~(~n_352 & n_3312);
 assign sub_485_2_n_1 = ~(n_373 & sub_485_2_n_28);
 assign sub_485_2_n_0 = ~(~n_657 & n_3319);
 assign n_1805 = (sub_504_2_n_74 ^ sub_504_2_n_147);
 assign n_1801 = ~(sub_504_2_n_102 | sub_504_2_n_148);
 assign n_1802 = ~(sub_504_2_n_77 ^ n_3575);
 assign n_1803 = ~(sub_504_2_n_17 ^ n_3576);
 assign sub_504_2_n_148 = ~(~sub_504_2_n_97 | sub_504_2_n_143);
 assign sub_504_2_n_147 = (~sub_504_2_n_54 | (n_3577 & sub_504_2_n_40));
 assign n_1806 = ~(n_3577 ^ sub_504_2_n_72);
 assign n_1807 = ~(sub_504_2_n_18 ^ n_3578);
 assign n_1809 = (sub_504_2_n_63 ^ n_3579);
 assign sub_504_2_n_143 = ~(sub_504_2_n_129 & (~sub_504_2_n_81 & ~sub_504_2_n_68));
 assign n_1804 = ~(sub_504_2_n_76 ^ sub_504_2_n_129);
 assign n_1808 = ~(sub_504_2_n_64 ^ sub_504_2_n_128);
 assign n_1810 = ~(sub_504_2_n_62 ^ n_3574);
 assign n_1811 = ~(sub_504_2_n_16 ^ n_3580);
 assign sub_504_2_n_129 = ~(~sub_504_2_n_106 & sub_504_2_n_127);
 assign sub_504_2_n_128 = ~(~sub_504_2_n_95 & sub_504_2_n_123);
 assign sub_504_2_n_127 = ~(sub_504_2_n_120 & (~sub_504_2_n_91 & ~sub_504_2_n_90));
 assign n_1812 = ~(sub_504_2_n_13 ^ sub_504_2_n_121);
 assign n_1813 = ~(sub_504_2_n_15 ^ n_3581);
 assign sub_504_2_n_123 = ~(~sub_504_2_n_90 & sub_504_2_n_121);
 assign sub_504_2_n_120 = ~(sub_504_2_n_115 & (~sub_504_2_n_46 & ~sub_504_2_n_93));
 assign sub_504_2_n_121 = ~(sub_504_2_n_115 & (~sub_504_2_n_46 & ~sub_504_2_n_93));
 assign n_1814 = ~(sub_504_2_n_75 ^ n_3582);
 assign n_1815 = ~(sub_504_2_n_19 ^ n_3583);
 assign sub_504_2_n_115 = ~(sub_504_2_n_109 & (~sub_504_2_n_70 & ~sub_504_2_n_84));
 assign n_1816 = ~(sub_504_2_n_61 ^ sub_504_2_n_109);
 assign sub_504_2_n_109 = ~(sub_504_2_n_107 & sub_504_2_n_60);
 assign n_1817 = (sub_504_2_n_20 ^ n_3584);
 assign sub_504_2_n_107 = ~(sub_504_2_n_59 & (sub_504_2_n_1 | (sub_504_2_n_101 & sub_504_2_n_51)));
 assign sub_504_2_n_106 = ~(sub_504_2_n_98 & (~sub_504_2_n_11 & ~sub_504_2_n_22));
 assign n_1818 = (sub_504_2_n_101 ^ sub_504_2_n_73);
 assign sub_504_2_n_102 = ~(sub_504_2_n_99 | n_3585);
 assign sub_504_2_n_101 = ((sub_485_2_n_27 & n_381) | (n_3058 & (sub_485_2_n_27 ^ n_381)));
 assign n_1819 = (n_3058 ^ (sub_485_2_n_27 ^ n_381));
 assign sub_504_2_n_99 = ~(~sub_504_2_n_68 & sub_504_2_n_96);
 assign sub_504_2_n_98 = ~(~sub_504_2_n_91 & sub_504_2_n_95);
 assign sub_504_2_n_97 = ~(~sub_504_2_n_96 | sub_504_2_n_67);
 assign sub_504_2_n_96 = ~(n_667 | (n_545 | (~sub_504_2_n_65 | ~sub_504_2_n_48)));
 assign sub_504_2_n_95 = ~(sub_504_2_n_89 & (~sub_504_2_n_82 | sub_504_2_n_88));
 assign sub_504_2_n_93 = ~(sub_504_2_n_78 & (sub_504_2_n_86 | sub_504_2_n_70));
 assign sub_504_2_n_91 = ~(sub_504_2_n_83 & sub_504_2_n_69);
 assign sub_504_2_n_90 = ~(sub_504_2_n_71 & sub_504_2_n_82);
 assign sub_504_2_n_89 = (~sub_504_2_n_4 & (sub_504_2_n_38 | sub_504_2_n_49));
 assign sub_504_2_n_88 = (~sub_504_2_n_10 & (sub_504_2_n_34 | sub_504_2_n_35));
 assign sub_504_2_n_86 = (~sub_504_2_n_2 & (sub_504_2_n_7 | sub_504_2_n_41));
 assign sub_504_2_n_78 = ~(sub_504_2_n_43 & sub_504_2_n_58);
 assign sub_504_2_n_84 = ~(sub_504_2_n_5 & sub_504_2_n_42);
 assign sub_504_2_n_77 = ~(sub_504_2_n_47 & sub_504_2_n_3);
 assign sub_504_2_n_83 = ~(sub_504_2_n_36 | sub_504_2_n_53);
 assign sub_504_2_n_76 = ~(sub_504_2_n_55 & sub_504_2_n_9);
 assign sub_504_2_n_75 = ~(sub_504_2_n_44 & sub_504_2_n_45);
 assign sub_504_2_n_74 = ~(sub_504_2_n_11 | sub_504_2_n_33);
 assign sub_504_2_n_73 = ~(sub_504_2_n_1 | sub_504_2_n_50);
 assign sub_504_2_n_72 = ~(sub_504_2_n_54 & sub_504_2_n_40);
 assign sub_504_2_n_82 = ~(sub_504_2_n_30 | sub_504_2_n_49);
 assign sub_504_2_n_81 = ~(~n_453 & sub_504_2_n_3);
 assign n_1820 = ~(sub_504_2_n_29 & (~{in2[13]} | {in1[0]}));
 assign sub_504_2_n_65 = ~(n_625 | (n_591 | (n_412 | n_504)));
 assign sub_504_2_n_64 = ~(sub_504_2_n_52 & sub_504_2_n_37);
 assign sub_504_2_n_63 = ~(sub_504_2_n_4 | sub_504_2_n_49);
 assign sub_504_2_n_62 = ~(sub_504_2_n_38 & sub_504_2_n_31);
 assign sub_504_2_n_71 = ~(sub_504_2_n_32 | sub_504_2_n_35);
 assign sub_504_2_n_70 = ~(sub_504_2_n_45 & sub_504_2_n_58);
 assign sub_504_2_n_69 = ~(sub_504_2_n_39 | sub_504_2_n_33);
 assign sub_504_2_n_61 = ~(sub_504_2_n_7 & sub_504_2_n_5);
 assign sub_504_2_n_68 = (n_483 | (n_601 | (n_341 | n_463)));
 assign sub_504_2_n_67 = ~(sub_504_2_n_9 & sub_504_2_n_57);
 assign sub_504_2_n_59 = ~sub_504_2_n_12;
 assign sub_504_2_n_57 = ~sub_504_2_n_56;
 assign sub_504_2_n_54 = ~sub_504_2_n_6;
 assign sub_504_2_n_51 = ~sub_504_2_n_50;
 assign sub_504_2_n_48 = ~(n_1112 | n_555);
 assign sub_504_2_n_60 = ~(~n_535 & n_3323);
 assign sub_504_2_n_58 = ~(sub_504_2_n_28 & n_680);
 assign sub_504_2_n_56 = ~(~n_565 | n_3327);
 assign sub_504_2_n_55 = ~(~n_473 & n_3328);
 assign sub_504_2_n_53 = ~(~n_352 | n_1788);
 assign sub_504_2_n_52 = ~(~n_690 & n_3732);
 assign sub_504_2_n_50 = ~(~n_422 | n_1799);
 assign sub_504_2_n_49 = ~(~n_432 | n_3733);
 assign sub_504_2_n_44 = ~sub_504_2_n_43;
 assign sub_504_2_n_42 = ~sub_504_2_n_41;
 assign sub_504_2_n_40 = ~sub_504_2_n_39;
 assign sub_504_2_n_37 = ~sub_504_2_n_36;
 assign sub_504_2_n_31 = ~sub_504_2_n_30;
 assign sub_504_2_n_47 = ~(~n_611 & n_1783);
 assign sub_504_2_n_46 = ~(n_680 | sub_504_2_n_28);
 assign sub_504_2_n_45 = ~(sub_504_2_n_26 & n_657);
 assign sub_504_2_n_43 = ~(n_657 | sub_504_2_n_26);
 assign sub_504_2_n_41 = ~(~n_639 | n_3322);
 assign sub_504_2_n_39 = ~(~n_373 | n_3324);
 assign sub_504_2_n_38 = ~(~n_362 & n_1791);
 assign sub_504_2_n_36 = ~(~n_690 | n_3732);
 assign sub_504_2_n_35 = ~(~n_398 | n_3326);
 assign sub_504_2_n_34 = ~(~n_442 & n_3329);
 assign sub_504_2_n_33 = ~(~n_524 | n_3321);
 assign sub_504_2_n_32 = ~(~n_442 | n_3329);
 assign sub_504_2_n_30 = ~(~n_362 | n_1791);
 assign sub_504_2_n_29 = ~({in1[0]} & ~{in2[13]});
 assign sub_504_2_n_28 = ~n_3330;
 assign sub_504_2_n_26 = ~n_3325;
 assign sub_504_2_n_22 = ~(sub_504_2_n_14 & (~sub_504_2_n_69 | n_3587));
 assign sub_504_2_n_20 = ~(~sub_504_2_n_60 | sub_504_2_n_12);
 assign sub_504_2_n_19 = ~(~sub_504_2_n_2 & sub_504_2_n_42);
 assign sub_504_2_n_18 = ~(sub_504_2_n_0 & ~sub_504_2_n_53);
 assign sub_504_2_n_17 = ~(~sub_504_2_n_8 & sub_504_2_n_57);
 assign sub_504_2_n_16 = (sub_504_2_n_10 | sub_504_2_n_35);
 assign sub_504_2_n_15 = ~(~sub_504_2_n_46 & sub_504_2_n_58);
 assign sub_504_2_n_14 = ~(sub_504_2_n_6 & ~sub_504_2_n_33);
 assign sub_504_2_n_13 = ~(sub_504_2_n_34 & ~sub_504_2_n_32);
 assign sub_504_2_n_12 = ~(n_3323 | ~n_535);
 assign sub_504_2_n_11 = ~(n_524 | ~n_3321);
 assign sub_504_2_n_10 = ~(n_398 | ~n_3326);
 assign sub_504_2_n_9 = ~(~n_3328 & n_473);
 assign sub_504_2_n_8 = ~(n_565 | ~n_3327);
 assign sub_504_2_n_7 = ~(~n_702 & n_3734);
 assign sub_504_2_n_6 = ~(n_373 | ~n_3324);
 assign sub_504_2_n_5 = ~(~n_3734 & n_702);
 assign sub_504_2_n_4 = ~(n_432 | ~n_3733);
 assign sub_504_2_n_3 = ~(~n_1783 & n_611);
 assign sub_504_2_n_2 = ~(n_639 | ~n_3322);
 assign sub_504_2_n_1 = ~(n_422 | ~n_1799);
 assign sub_504_2_n_0 = ~(~n_352 & n_1788);
 assign sub_523_2_n_27 = (~sub_523_2_n_94 | (sub_523_2_n_74 & sub_523_2_n_131));
 assign n_1841 = ~(sub_523_2_n_82 ^ n_3588);
 assign n_1845 = (sub_523_2_n_21 ^ sub_523_2_n_17);
 assign n_1842 = ~(sub_523_2_n_81 ^ sub_523_2_n_27);
 assign n_1843 = ~(sub_523_2_n_23 ^ n_3589);
 assign n_1846 = ~(sub_523_2_n_139 ^ sub_523_2_n_78);
 assign n_1847 = (sub_523_2_n_20 ^ n_3591);
 assign n_1849 = ~(sub_523_2_n_16 ^ sub_523_2_n_136);
 assign n_1844 = ~(sub_523_2_n_79 ^ sub_523_2_n_131);
 assign sub_523_2_n_139 = ~(sub_523_2_n_92 & (~sub_523_2_n_86 | n_3592));
 assign sub_523_2_n_136 = ~(sub_523_2_n_11 & (sub_523_2_n_24 | sub_523_2_n_55));
 assign n_1848 = ~(n_3592 ^ sub_523_2_n_68);
 assign n_1850 = (sub_523_2_n_19 ^ sub_523_2_n_24);
 assign n_1851 = ~(sub_523_2_n_13 ^ sub_523_2_n_128);
 assign sub_523_2_n_131 = ~(sub_523_2_n_129 & sub_523_2_n_111);
 assign sub_523_2_n_129 = ~(sub_523_2_n_124 & (~sub_523_2_n_95 & ~sub_523_2_n_96));
 assign sub_523_2_n_128 = ~(sub_523_2_n_39 & (sub_523_2_n_123 | sub_523_2_n_38));
 assign n_1852 = (sub_523_2_n_14 ^ sub_523_2_n_123);
 assign n_1853 = ~(sub_523_2_n_18 ^ n_3593);
 assign sub_523_2_n_123 = ~sub_523_2_n_124;
 assign sub_523_2_n_124 = ~(sub_523_2_n_118 & (~sub_523_2_n_50 & ~sub_523_2_n_100));
 assign n_1854 = (sub_523_2_n_80 ^ n_3596);
 assign n_1855 = (sub_523_2_n_69 ^ sub_523_2_n_26);
 assign sub_523_2_n_118 = ~(n_3701 & (~sub_523_2_n_76 & ~sub_523_2_n_22));
 assign n_1856 = ~(sub_523_2_n_67 ^ n_3701);
 assign n_1857 = (sub_523_2_n_83 ^ n_3594);
 assign sub_523_2_n_112 = ~(sub_523_2_n_103 | (~sub_523_2_n_75 | ~sub_523_2_n_102));
 assign sub_523_2_n_111 = ~(sub_523_2_n_105 | (~sub_523_2_n_64 | ~n_3595));
 assign n_1858 = (n_840 ^ sub_523_2_n_15);
 assign sub_523_2_n_107 = ((sub_485_2_n_27 & n_402) | (n_3059 & (sub_485_2_n_27 ^ n_402)));
 assign n_1859 = (n_3059 ^ (sub_485_2_n_27 ^ n_402));
 assign sub_523_2_n_105 = ~(sub_523_2_n_101 | sub_523_2_n_96);
 assign sub_523_2_n_103 = ~(sub_523_2_n_98 | (~sub_523_2_n_71 | ~sub_523_2_n_4));
 assign sub_523_2_n_102 = ~(n_666 | (n_544 | (~n_3147 | ~n_3146)));
 assign sub_523_2_n_101 = ~(sub_523_2_n_93 | (sub_523_2_n_90 & sub_523_2_n_85));
 assign sub_523_2_n_100 = ~(sub_523_2_n_84 & (sub_523_2_n_89 | sub_523_2_n_76));
 assign sub_523_2_n_98 = ~(~sub_523_2_n_87 | sub_523_2_n_94);
 assign sub_523_2_n_96 = ~(sub_523_2_n_86 & sub_523_2_n_88);
 assign sub_523_2_n_95 = ~(sub_523_2_n_77 & sub_523_2_n_85);
 assign sub_523_2_n_94 = (~sub_523_2_n_10 & (sub_523_2_n_49 | sub_523_2_n_45));
 assign sub_523_2_n_93 = ~(sub_523_2_n_7 & (sub_523_2_n_11 | sub_523_2_n_42));
 assign sub_523_2_n_92 = ~sub_523_2_n_91;
 assign sub_523_2_n_91 = ~(sub_523_2_n_1 & (sub_523_2_n_12 | sub_523_2_n_60));
 assign sub_523_2_n_90 = ~(sub_523_2_n_2 & (sub_523_2_n_39 | sub_523_2_n_35));
 assign sub_523_2_n_89 = (~sub_523_2_n_8 & (sub_523_2_n_5 | sub_523_2_n_63));
 assign sub_523_2_n_84 = ~(sub_523_2_n_47 & sub_523_2_n_48);
 assign sub_523_2_n_88 = ~(sub_523_2_n_58 | sub_523_2_n_62);
 assign sub_523_2_n_87 = ~(sub_523_2_n_56 | sub_523_2_n_33);
 assign sub_523_2_n_83 = ~(sub_523_2_n_6 | sub_523_2_n_65);
 assign sub_523_2_n_82 = ~(sub_523_2_n_4 & sub_523_2_n_34);
 assign sub_523_2_n_86 = ~(sub_523_2_n_53 | sub_523_2_n_60);
 assign sub_523_2_n_81 = ~(sub_523_2_n_40 & sub_523_2_n_57);
 assign sub_523_2_n_80 = ~(sub_523_2_n_47 | sub_523_2_n_36);
 assign sub_523_2_n_79 = ~(sub_523_2_n_49 & sub_523_2_n_44);
 assign sub_523_2_n_85 = ~(sub_523_2_n_55 | sub_523_2_n_42);
 assign sub_523_2_n_78 = ~(sub_523_2_n_0 & sub_523_2_n_59);
 assign n_1860 = ~(sub_523_2_n_52 & (~{in2[12]} | {in1[0]}));
 assign sub_523_2_n_71 = ~(sub_523_2_n_9 & sub_523_2_n_34);
 assign sub_523_2_n_69 = ~(sub_523_2_n_8 | sub_523_2_n_63);
 assign sub_523_2_n_77 = ~(sub_523_2_n_38 | sub_523_2_n_35);
 assign sub_523_2_n_76 = ~(sub_523_2_n_37 & sub_523_2_n_48);
 assign sub_523_2_n_68 = ~(sub_523_2_n_61 | sub_523_2_n_53);
 assign sub_523_2_n_75 = ~(n_482 | (n_600 | (n_340 | n_462)));
 assign sub_523_2_n_67 = ~(sub_523_2_n_5 & sub_523_2_n_3);
 assign sub_523_2_n_74 = ~(sub_523_2_n_43 | sub_523_2_n_45);
 assign sub_523_2_n_61 = ~sub_523_2_n_12;
 assign sub_523_2_n_59 = ~sub_523_2_n_58;
 assign sub_523_2_n_57 = ~sub_523_2_n_56;
 assign sub_523_2_n_65 = ~(~n_534 | n_841);
 assign sub_523_2_n_64 = ~(~n_523 & n_850);
 assign sub_523_2_n_63 = ~(~n_638 | n_838);
 assign sub_523_2_n_62 = ~(~n_523 | n_850);
 assign sub_523_2_n_60 = ~(~n_351 | n_836);
 assign sub_523_2_n_58 = ~(~n_372 | n_848);
 assign sub_523_2_n_56 = ~(~n_610 | n_851);
 assign sub_523_2_n_55 = ~(~n_361 | n_834);
 assign sub_523_2_n_54 = ~(n_421 | sub_523_2_n_32);
 assign sub_523_2_n_53 = ~(~n_689 | n_835);
 assign sub_523_2_n_52 = ~({in1[0]} & ~{in2[12]});
 assign sub_523_2_n_47 = ~sub_523_2_n_46;
 assign sub_523_2_n_44 = ~sub_523_2_n_43;
 assign sub_523_2_n_40 = ~sub_523_2_n_9;
 assign sub_523_2_n_37 = ~sub_523_2_n_36;
 assign sub_523_2_n_34 = ~sub_523_2_n_33;
 assign sub_523_2_n_50 = ~(n_679 | sub_523_2_n_29);
 assign sub_523_2_n_49 = ~(~n_472 & n_846);
 assign sub_523_2_n_48 = ~(sub_523_2_n_29 & n_679);
 assign sub_523_2_n_46 = ~(~n_656 & n_845);
 assign sub_523_2_n_45 = ~(~n_564 | n_853);
 assign sub_523_2_n_43 = ~(~n_472 | n_846);
 assign sub_523_2_n_42 = ~(~n_431 | n_833);
 assign sub_523_2_n_41 = ~(sub_523_2_n_32 & n_421);
 assign sub_523_2_n_39 = ~(sub_523_2_n_31 & n_847);
 assign sub_523_2_n_38 = ~(n_847 | sub_523_2_n_31);
 assign sub_523_2_n_36 = ~(~n_656 | n_845);
 assign sub_523_2_n_35 = ~(~n_397 | n_837);
 assign sub_523_2_n_33 = ~(~n_452 | n_849);
 assign sub_523_2_n_32 = ~n_842;
 assign sub_523_2_n_31 = ~n_441;
 assign sub_523_2_n_29 = ~n_844;
 assign sub_523_2_n_26 = (~sub_523_2_n_5 | (sub_523_2_n_3 & n_3701));
 assign sub_523_2_n_24 = ~(sub_523_2_n_90 | (sub_523_2_n_77 & sub_523_2_n_124));
 assign sub_523_2_n_23 = (sub_523_2_n_10 | sub_523_2_n_45);
 assign sub_523_2_n_22 = ~(sub_523_2_n_3 & ~sub_523_2_n_63);
 assign sub_523_2_n_21 = ~(sub_523_2_n_64 & ~sub_523_2_n_62);
 assign sub_523_2_n_20 = ~(sub_523_2_n_1 & ~sub_523_2_n_60);
 assign sub_523_2_n_19 = ~(sub_523_2_n_11 & ~sub_523_2_n_55);
 assign sub_523_2_n_18 = ~(~sub_523_2_n_50 & sub_523_2_n_48);
 assign sub_523_2_n_17 = (sub_523_2_n_0 & ~(sub_523_2_n_139 & sub_523_2_n_59));
 assign sub_523_2_n_16 = ~(sub_523_2_n_7 & ~sub_523_2_n_42);
 assign sub_523_2_n_15 = ~(sub_523_2_n_54 | ~sub_523_2_n_41);
 assign sub_523_2_n_14 = ~(sub_523_2_n_39 & ~sub_523_2_n_38);
 assign sub_523_2_n_13 = ~(sub_523_2_n_2 & ~sub_523_2_n_35);
 assign sub_523_2_n_12 = ~(~n_689 & n_835);
 assign sub_523_2_n_11 = ~(~n_361 & n_834);
 assign sub_523_2_n_10 = ~(n_564 | ~n_853);
 assign sub_523_2_n_9 = ~(n_610 | ~n_851);
 assign sub_523_2_n_8 = ~(n_638 | ~n_838);
 assign sub_523_2_n_7 = ~(~n_431 & n_833);
 assign sub_523_2_n_6 = ~(n_534 | ~n_841);
 assign sub_523_2_n_5 = ~(~n_701 & n_852);
 assign sub_523_2_n_4 = ~(~n_452 & n_849);
 assign sub_523_2_n_3 = ~(~n_852 & n_701);
 assign sub_523_2_n_2 = ~(~n_397 & n_837);
 assign sub_523_2_n_1 = ~(~n_351 & n_836);
 assign sub_523_2_n_0 = ~(~n_372 & n_848);
 assign n_1896 = ~(sub_542_2_n_14 ^ sub_542_2_n_125);
 assign n_1883 = (sub_542_2_n_87 ^ sub_542_2_n_162);
 assign n_1887 = ~(sub_542_2_n_15 ^ n_3608);
 assign sub_542_2_n_162 = (~sub_542_2_n_54 | (sub_542_2_n_25 & sub_542_2_n_8));
 assign n_1882 = ~(sub_542_2_n_88 ^ sub_542_2_n_28);
 assign n_1884 = ~(sub_542_2_n_86 ^ sub_542_2_n_25);
 assign n_1885 = ~(sub_542_2_n_23 ^ n_3597);
 assign n_1888 = (sub_542_2_n_78 ^ n_3599);
 assign n_1889 = ~(sub_542_2_n_77 ^ n_3598);
 assign n_1891 = ~(sub_542_2_n_16 ^ n_3601);
 assign n_1881 = ~(sub_542_2_n_118 | n_3600);
 assign n_1892 = ~(sub_542_2_n_74 ^ sub_542_2_n_137);
 assign n_1890 = ~(sub_542_2_n_76 ^ n_3602);
 assign n_1886 = ~(sub_542_2_n_85 ^ sub_542_2_n_135);
 assign n_1893 = ~(sub_542_2_n_75 ^ n_3603);
 assign sub_542_2_n_137 = ~(~sub_542_2_n_100 & sub_542_2_n_132);
 assign sub_542_2_n_135 = ~(sub_542_2_n_116 & n_3604);
 assign n_1894 = ~(sub_542_2_n_73 ^ sub_542_2_n_129);
 assign n_1895 = (sub_542_2_n_21 ^ sub_542_2_n_128);
 assign sub_542_2_n_132 = ~(~sub_542_2_n_82 & sub_542_2_n_129);
 assign sub_542_2_n_129 = ~(sub_542_2_n_126 & (~sub_542_2_n_48 & ~sub_542_2_n_107));
 assign sub_542_2_n_128 = ~(sub_542_2_n_38 & (~sub_542_2_n_39 | sub_542_2_n_125));
 assign n_1897 = ~(sub_542_2_n_71 ^ n_3605);
 assign sub_542_2_n_126 = ~(n_3703 & (~sub_542_2_n_92 & ~sub_542_2_n_83));
 assign sub_542_2_n_125 = ~(sub_542_2_n_101 | (~sub_542_2_n_92 & n_3703));
 assign n_1898 = (sub_542_2_n_18 ^ n_3703);
 assign n_1899 = (sub_542_2_n_72 ^ n_3606);
 assign sub_542_2_n_118 = ~(sub_542_2_n_110 | (sub_542_2_n_111 & sub_542_2_n_22));
 assign sub_542_2_n_116 = ~(sub_542_2_n_49 | (sub_542_2_n_108 | (sub_542_2_n_24 & sub_542_2_n_104)));
 assign n_1900 = (sub_542_2_n_113 ^ sub_542_2_n_84);
 assign sub_542_2_n_113 = ((sub_561_2_n_34 & n_495) | (n_3358 & (sub_561_2_n_34 ^ n_495)));
 assign n_1901 = (n_3358 ^ (sub_561_2_n_34 ^ n_495));
 assign sub_542_2_n_111 = ~(~sub_542_2_n_102 & sub_542_2_n_109);
 assign sub_542_2_n_110 = ~(n_3147 & (n_3146 & (~n_666 & ~n_544)));
 assign sub_542_2_n_109 = ~(sub_542_2_n_97 & (sub_542_2_n_99 | sub_542_2_n_19));
 assign sub_542_2_n_108 = ~(sub_542_2_n_79 & (n_3607 | sub_542_2_n_95));
 assign sub_542_2_n_107 = ~(sub_542_2_n_89 & (sub_542_2_n_17 | sub_542_2_n_83));
 assign sub_542_2_n_104 = ~(sub_542_2_n_94 | sub_542_2_n_95);
 assign sub_542_2_n_103 = ~(sub_542_2_n_82 | sub_542_2_n_91);
 assign sub_542_2_n_102 = ~(~n_600 & (n_3148 & sub_542_2_n_1));
 assign sub_542_2_n_101 = ~sub_542_2_n_17;
 assign sub_542_2_n_97 = (~sub_542_2_n_10 & (sub_542_2_n_54 | sub_542_2_n_60));
 assign sub_542_2_n_96 = (~sub_542_2_n_9 & (sub_542_2_n_53 | sub_542_2_n_44));
 assign sub_542_2_n_100 = ~(sub_542_2_n_50 & (sub_542_2_n_42 | sub_542_2_n_45));
 assign sub_542_2_n_99 = (~sub_542_2_n_7 & (sub_542_2_n_47 | sub_542_2_n_35));
 assign sub_542_2_n_89 = ~(sub_542_2_n_37 & sub_542_2_n_65);
 assign sub_542_2_n_95 = ~(sub_542_2_n_64 & sub_542_2_n_59);
 assign sub_542_2_n_88 = ~(sub_542_2_n_66 & sub_542_2_n_1);
 assign sub_542_2_n_94 = ~(sub_542_2_n_13 & sub_542_2_n_56);
 assign sub_542_2_n_87 = ~(sub_542_2_n_10 | sub_542_2_n_60);
 assign sub_542_2_n_93 = ~(sub_542_2_n_0 & sub_542_2_n_36);
 assign sub_542_2_n_86 = ~(sub_542_2_n_54 & sub_542_2_n_8);
 assign sub_542_2_n_92 = ~(sub_542_2_n_58 & sub_542_2_n_41);
 assign sub_542_2_n_85 = ~(sub_542_2_n_47 & sub_542_2_n_0);
 assign sub_542_2_n_91 = ~(~sub_542_2_n_44 & sub_542_2_n_4);
 assign sub_542_2_n_84 = ~(sub_542_2_n_6 | sub_542_2_n_61);
 assign n_1902 = ~(sub_542_2_n_52 & (~{in2[11]} | {in1[0]}));
 assign sub_542_2_n_79 = ~(sub_542_2_n_11 & sub_542_2_n_59);
 assign sub_542_2_n_78 = ~(sub_542_2_n_11 | sub_542_2_n_63);
 assign sub_542_2_n_77 = ~(sub_542_2_n_67 & sub_542_2_n_56);
 assign sub_542_2_n_83 = ~(sub_542_2_n_39 & sub_542_2_n_65);
 assign sub_542_2_n_76 = ~(sub_542_2_n_43 & sub_542_2_n_13);
 assign sub_542_2_n_75 = ~(sub_542_2_n_50 & sub_542_2_n_46);
 assign sub_542_2_n_74 = ~(sub_542_2_n_53 & sub_542_2_n_4);
 assign sub_542_2_n_82 = ~(sub_542_2_n_2 & sub_542_2_n_46);
 assign sub_542_2_n_73 = ~(sub_542_2_n_42 & sub_542_2_n_2);
 assign sub_542_2_n_72 = ~(sub_542_2_n_12 | sub_542_2_n_69);
 assign sub_542_2_n_71 = ~(sub_542_2_n_5 & sub_542_2_n_41);
 assign sub_542_2_n_64 = ~sub_542_2_n_63;
 assign sub_542_2_n_62 = ~sub_542_2_n_61;
 assign sub_542_2_n_58 = ~sub_542_2_n_57;
 assign sub_542_2_n_56 = ~sub_542_2_n_55;
 assign sub_542_2_n_69 = ~(~n_534 | n_3353);
 assign sub_542_2_n_67 = ~(~n_351 & n_3347);
 assign sub_542_2_n_66 = ~(~n_482 & n_3343);
 assign sub_542_2_n_65 = ~(sub_542_2_n_33 & n_679);
 assign sub_542_2_n_63 = ~(~n_372 | n_3345);
 assign sub_542_2_n_61 = ~(~n_421 | n_3355);
 assign sub_542_2_n_60 = ~(~n_452 | n_3356);
 assign sub_542_2_n_59 = ~(sub_542_2_n_31 & n_523);
 assign sub_542_2_n_57 = ~(~n_701 | n_3352);
 assign sub_542_2_n_55 = ~(~n_351 | n_3347);
 assign sub_542_2_n_54 = ~(~n_610 & n_3357);
 assign sub_542_2_n_53 = ~(~n_361 & n_3360);
 assign sub_542_2_n_52 = ~({in1[0]} & ~{in2[11]});
 assign sub_542_2_n_46 = ~sub_542_2_n_45;
 assign sub_542_2_n_41 = ~sub_542_2_n_40;
 assign sub_542_2_n_38 = ~sub_542_2_n_37;
 assign sub_542_2_n_36 = ~sub_542_2_n_35;
 assign sub_542_2_n_50 = ~(~n_397 & n_3361);
 assign sub_542_2_n_49 = ~(n_523 | sub_542_2_n_31);
 assign sub_542_2_n_48 = ~(n_679 | sub_542_2_n_33);
 assign sub_542_2_n_47 = ~(~n_472 & n_3350);
 assign sub_542_2_n_45 = ~(~n_397 | n_3361);
 assign sub_542_2_n_44 = ~(~n_431 | n_3354);
 assign sub_542_2_n_43 = ~(~n_689 & n_3351);
 assign sub_542_2_n_42 = ~(~n_441 & n_3362);
 assign sub_542_2_n_40 = ~(~n_638 | n_3349);
 assign sub_542_2_n_39 = ~(sub_542_2_n_34 & n_656);
 assign sub_542_2_n_37 = ~(n_656 | sub_542_2_n_34);
 assign sub_542_2_n_35 = ~(~n_564 | n_3344);
 assign sub_542_2_n_34 = ~n_3348;
 assign sub_542_2_n_33 = ~n_3346;
 assign sub_542_2_n_31 = ~n_3359;
 assign sub_542_2_n_28 = ~(n_3692 & ~sub_542_2_n_109);
 assign sub_542_2_n_25 = ~(sub_542_2_n_99 & (~sub_542_2_n_135 | sub_542_2_n_93));
 assign sub_542_2_n_24 = ~(sub_542_2_n_96 & (~sub_542_2_n_100 | sub_542_2_n_91));
 assign sub_542_2_n_23 = ~(~sub_542_2_n_7 & sub_542_2_n_36);
 assign sub_542_2_n_22 = ~(n_3148 & (~sub_542_2_n_66 & ~n_600));
 assign sub_542_2_n_21 = ~(sub_542_2_n_48 | ~sub_542_2_n_65);
 assign sub_542_2_n_19 = ~(sub_542_2_n_8 & ~sub_542_2_n_60);
 assign sub_542_2_n_18 = ~(~sub_542_2_n_3 | sub_542_2_n_57);
 assign sub_542_2_n_17 = (sub_542_2_n_5 & (sub_542_2_n_3 | sub_542_2_n_40));
 assign sub_542_2_n_16 = (sub_542_2_n_9 | sub_542_2_n_44);
 assign sub_542_2_n_15 = ~(~sub_542_2_n_49 & sub_542_2_n_59);
 assign sub_542_2_n_14 = ~(sub_542_2_n_37 | ~sub_542_2_n_39);
 assign sub_542_2_n_13 = ~(~n_3351 & n_689);
 assign sub_542_2_n_12 = ~(n_534 | ~n_3353);
 assign sub_542_2_n_11 = ~(n_372 | ~n_3345);
 assign sub_542_2_n_10 = ~(n_452 | ~n_3356);
 assign sub_542_2_n_9 = ~(n_431 | ~n_3354);
 assign sub_542_2_n_8 = ~(~n_3357 & n_610);
 assign sub_542_2_n_7 = ~(n_564 | ~n_3344);
 assign sub_542_2_n_6 = ~(n_421 | ~n_3355);
 assign sub_542_2_n_5 = ~(~n_638 & n_3349);
 assign sub_542_2_n_4 = ~(~n_3360 & n_361);
 assign sub_542_2_n_3 = ~(~n_701 & n_3352);
 assign sub_542_2_n_2 = ~(~n_3362 & n_441);
 assign sub_542_2_n_1 = ~(~n_3343 & n_482);
 assign sub_542_2_n_0 = ~(~n_3350 & n_472);
 assign n_1924 = ~(n_3152 & sub_561_2_n_172);
 assign n_1925 = ~(n_905 ^ n_3609);
 assign n_1927 = ~(n_890 ^ n_3610);
 assign sub_561_2_n_172 = ~(sub_561_2_n_163 | (~n_3150 | ~n_3149));
 assign n_1931 = (n_908 ^ sub_561_2_n_25);
 assign n_1926 = ~(sub_561_2_n_91 ^ n_3611);
 assign n_1928 = (n_886 ^ n_3612);
 assign n_1929 = ~(n_873 ^ n_3613);
 assign sub_561_2_n_163 = ~(n_904 | (n_903 & (n_893 & n_906)));
 assign n_1932 = (sub_561_2_n_153 ^ sub_561_2_n_78);
 assign n_1935 = ~(n_858 ^ n_898);
 assign n_1930 = ~(sub_561_2_n_87 ^ n_906);
 assign sub_561_2_n_153 = ~(n_897 & (n_894 | n_892));
 assign sub_561_2_n_152 = ~(sub_561_2_n_10 & (n_3212 | sub_561_2_n_44));
 assign n_1934 = (sub_561_2_n_76 ^ n_894);
 assign n_1936 = (sub_561_2_n_19 ^ n_3212);
 assign n_1937 = (sub_561_2_n_15 ^ sub_561_2_n_143);
 assign sub_561_2_n_145 = ~(sub_561_2_n_139 & (~sub_561_2_n_111 & ~sub_561_2_n_109));
 assign sub_561_2_n_143 = ~(sub_561_2_n_52 | (~sub_561_2_n_43 & sub_561_2_n_139));
 assign n_1938 = (sub_561_2_n_18 ^ sub_561_2_n_138);
 assign n_1939 = (sub_561_2_n_74 ^ sub_561_2_n_137);
 assign sub_561_2_n_138 = ~sub_561_2_n_139;
 assign sub_561_2_n_139 = ~(sub_561_2_n_133 & (~sub_561_2_n_13 & ~sub_561_2_n_115));
 assign sub_561_2_n_137 = ~(sub_561_2_n_60 & (~sub_561_2_n_36 | sub_561_2_n_132));
 assign n_1941 = ~(sub_561_2_n_77 ^ n_3616);
 assign n_1940 = (sub_561_2_n_75 ^ sub_561_2_n_132);
 assign sub_561_2_n_133 = ~(n_3707 & (~sub_561_2_n_97 & ~sub_561_2_n_99));
 assign sub_561_2_n_132 = ~(sub_561_2_n_107 | (~sub_561_2_n_99 & n_3707));
 assign n_1942 = ~(sub_561_2_n_88 ^ n_3707);
 assign n_1943 = (sub_561_2_n_90 ^ n_3617);
 assign n_1944 = (sub_561_2_n_121 ^ sub_561_2_n_89);
 assign sub_561_2_n_122 = ~(sub_561_2_n_113 & (n_3618 | sub_561_2_n_21));
 assign sub_561_2_n_121 = ((sub_561_2_n_34 & n_709) | (n_3377 & (sub_561_2_n_34 ^ n_709)));
 assign n_1945 = (n_3377 ^ (sub_561_2_n_34 ^ n_709));
 assign sub_561_2_n_119 = ~(sub_561_2_n_117 | sub_561_2_n_111);
 assign sub_561_2_n_117 = ~(sub_561_2_n_101 | (sub_561_2_n_104 & sub_561_2_n_85));
 assign sub_561_2_n_115 = ~(sub_561_2_n_80 & (sub_561_2_n_26 | sub_561_2_n_97));
 assign sub_561_2_n_113 = ~(sub_561_2_n_102 & n_3148);
 assign sub_561_2_n_110 = ~sub_561_2_n_21;
 assign sub_561_2_n_112 = ~(sub_561_2_n_86 | sub_561_2_n_100);
 assign sub_561_2_n_111 = ~(sub_561_2_n_95 & sub_561_2_n_98);
 assign sub_561_2_n_109 = ~(sub_561_2_n_83 & sub_561_2_n_85);
 assign sub_561_2_n_107 = ~sub_561_2_n_26;
 assign sub_561_2_n_106 = ~sub_561_2_n_105;
 assign sub_561_2_n_102 = ~(sub_561_2_n_5 & (sub_561_2_n_42 | sub_561_2_n_38));
 assign sub_561_2_n_101 = ~(sub_561_2_n_8 & (sub_561_2_n_10 | sub_561_2_n_49));
 assign sub_561_2_n_105 = ~(sub_561_2_n_3 & (sub_561_2_n_4 | sub_561_2_n_56));
 assign sub_561_2_n_104 = ~(sub_561_2_n_12 & (sub_561_2_n_7 | sub_561_2_n_37));
 assign sub_561_2_n_96 = ~sub_561_2_n_95;
 assign sub_561_2_n_100 = ~(sub_561_2_n_58 & sub_561_2_n_51);
 assign sub_561_2_n_92 = ~(sub_561_2_n_70 & sub_561_2_n_51);
 assign sub_561_2_n_99 = ~(sub_561_2_n_6 & sub_561_2_n_46);
 assign sub_561_2_n_98 = ~(sub_561_2_n_67 | sub_561_2_n_40);
 assign sub_561_2_n_97 = ~(sub_561_2_n_36 & sub_561_2_n_48);
 assign sub_561_2_n_95 = ~(sub_561_2_n_64 | sub_561_2_n_56);
 assign sub_561_2_n_91 = ~(n_862 & n_863);
 assign sub_561_2_n_90 = ~(sub_561_2_n_1 | sub_561_2_n_68);
 assign sub_561_2_n_89 = ~(sub_561_2_n_11 | sub_561_2_n_61);
 assign sub_561_2_n_88 = ~(sub_561_2_n_2 & sub_561_2_n_6);
 assign sub_561_2_n_87 = ~(n_857 & n_859);
 assign n_1946 = ~(sub_561_2_n_55 & (~{in2[10]} | {in1[0]}));
 assign sub_561_2_n_80 = ~(sub_561_2_n_59 & sub_561_2_n_48);
 assign sub_561_2_n_78 = ~(n_907 | n_910);
 assign sub_561_2_n_77 = ~(sub_561_2_n_71 & sub_561_2_n_46);
 assign sub_561_2_n_76 = ~(n_899 & n_895);
 assign sub_561_2_n_75 = ~(sub_561_2_n_60 & sub_561_2_n_36);
 assign sub_561_2_n_86 = ~(sub_561_2_n_9 & sub_561_2_n_41);
 assign sub_561_2_n_74 = ~(sub_561_2_n_13 | sub_561_2_n_47);
 assign sub_561_2_n_85 = ~(sub_561_2_n_44 | sub_561_2_n_49);
 assign sub_561_2_n_83 = ~(sub_561_2_n_43 | sub_561_2_n_37);
 assign sub_561_2_n_66 = ~sub_561_2_n_0;
 assign sub_561_2_n_65 = ~sub_561_2_n_64;
 assign sub_561_2_n_62 = ~sub_561_2_n_61;
 assign sub_561_2_n_60 = ~sub_561_2_n_59;
 assign sub_561_2_n_58 = ~sub_561_2_n_57;
 assign sub_561_2_n_73 = ~(n_564 | sub_561_2_n_32);
 assign sub_561_2_n_72 = ~(~n_523 & n_3365);
 assign sub_561_2_n_71 = ~(sub_561_2_n_31 & n_3371);
 assign sub_561_2_n_70 = ~(sub_561_2_n_30 & n_3375);
 assign sub_561_2_n_68 = ~(~n_534 | n_1921);
 assign sub_561_2_n_67 = ~(~n_372 | n_3366);
 assign sub_561_2_n_64 = ~(~n_689 | n_3373);
 assign sub_561_2_n_63 = ~(~n_610 & n_3364);
 assign sub_561_2_n_61 = ~(~n_421 | n_3372);
 assign sub_561_2_n_59 = ~(n_656 | sub_561_2_n_33);
 assign sub_561_2_n_57 = ~(~n_610 | n_3364);
 assign sub_561_2_n_56 = ~(~n_351 | n_3370);
 assign sub_561_2_n_55 = ~({in1[0]} & ~{in2[10]});
 assign sub_561_2_n_52 = ~sub_561_2_n_7;
 assign sub_561_2_n_51 = ~sub_561_2_n_50;
 assign sub_561_2_n_48 = ~sub_561_2_n_47;
 assign sub_561_2_n_46 = ~sub_561_2_n_45;
 assign sub_561_2_n_50 = ~(n_3375 | sub_561_2_n_30);
 assign sub_561_2_n_49 = ~(~n_431 | n_3379);
 assign sub_561_2_n_47 = ~(~n_679 | n_3367);
 assign sub_561_2_n_45 = ~(n_3371 | sub_561_2_n_31);
 assign sub_561_2_n_44 = ~(~n_361 | n_3380);
 assign sub_561_2_n_43 = ~(~n_441 | n_1916);
 assign sub_561_2_n_42 = ~(~n_482 & n_3374);
 assign sub_561_2_n_41 = ~(sub_561_2_n_32 & n_564);
 assign sub_561_2_n_40 = ~(~n_523 | n_3365);
 assign sub_561_2_n_39 = ~(~n_472 & n_3378);
 assign sub_561_2_n_38 = ~(~n_600 | n_3363);
 assign sub_561_2_n_37 = ~(~n_397 | n_3381);
 assign sub_561_2_n_36 = ~(sub_561_2_n_33 & n_656);
 assign sub_561_2_n_34 = ~n_387;
 assign sub_561_2_n_33 = ~n_3368;
 assign sub_561_2_n_32 = ~n_3369;
 assign sub_561_2_n_31 = ~n_638;
 assign sub_561_2_n_30 = ~n_452;
 assign sub_561_2_n_27 = ~(~sub_561_2_n_73 & sub_561_2_n_41);
 assign sub_561_2_n_26 = (sub_561_2_n_71 & (sub_561_2_n_2 | sub_561_2_n_45));
 assign sub_561_2_n_25 = ~(n_907 | (~n_910 & sub_561_2_n_153));
 assign sub_561_2_n_24 = ~(~sub_561_2_n_63 | sub_561_2_n_57);
 assign sub_561_2_n_22 = ~(sub_561_2_n_3 & ~sub_561_2_n_56);
 assign sub_561_2_n_21 = ~(sub_561_2_n_14 & (n_3148 & ~sub_561_2_n_38));
 assign sub_561_2_n_20 = ~(sub_561_2_n_8 & ~sub_561_2_n_49);
 assign sub_561_2_n_19 = ~(sub_561_2_n_10 & ~sub_561_2_n_44);
 assign sub_561_2_n_18 = ~(sub_561_2_n_7 & ~sub_561_2_n_43);
 assign sub_561_2_n_17 = ~(sub_561_2_n_72 & ~sub_561_2_n_40);
 assign sub_561_2_n_16 = ~(sub_561_2_n_5 & ~sub_561_2_n_38);
 assign sub_561_2_n_15 = ~(sub_561_2_n_12 & ~sub_561_2_n_37);
 assign sub_561_2_n_14 = ~(~n_3374 & n_482);
 assign sub_561_2_n_13 = ~(n_679 | ~n_3367);
 assign sub_561_2_n_12 = ~(~n_397 & n_3381);
 assign sub_561_2_n_11 = ~(n_421 | ~n_3372);
 assign sub_561_2_n_10 = ~(~n_361 & n_3380);
 assign sub_561_2_n_9 = ~(~n_3378 & n_472);
 assign sub_561_2_n_8 = ~(~n_431 & n_3379);
 assign sub_561_2_n_7 = ~(~n_441 & n_1916);
 assign sub_561_2_n_6 = ~(~n_3376 & n_701);
 assign sub_561_2_n_5 = ~(~n_600 & n_3363);
 assign sub_561_2_n_4 = ~(~n_689 & n_3373);
 assign sub_561_2_n_3 = ~(~n_351 & n_3370);
 assign sub_561_2_n_2 = ~(~n_701 & n_3376);
 assign sub_561_2_n_1 = ~(n_534 | ~n_1921);
 assign sub_561_2_n_0 = ~(~n_372 & n_3366);
 assign n_1986 = ~(sub_580_2_n_27 ^ sub_580_2_n_127);
 assign n_1969 = ~sub_580_2_n_174;
 assign sub_580_2_n_174 = ~(~n_3152 | sub_580_2_n_170);
 assign n_1970 = ~(sub_580_2_n_26 ^ n_3622);
 assign n_1971 = ~(sub_580_2_n_30 ^ n_3623);
 assign n_1973 = ~(sub_580_2_n_28 ^ n_3624);
 assign sub_580_2_n_170 = ~(sub_580_2_n_160 & (~sub_580_2_n_85 & ~sub_580_2_n_43));
 assign n_1977 = ~(sub_580_2_n_31 ^ n_3625);
 assign n_1972 = ~(sub_580_2_n_29 ^ sub_580_2_n_153);
 assign n_1974 = (sub_580_2_n_19 ^ n_3626);
 assign n_1975 = ~(sub_580_2_n_22 ^ n_3627);
 assign sub_580_2_n_160 = ~(sub_580_2_n_154 & sub_580_2_n_118);
 assign n_1978 = ~(sub_580_2_n_83 ^ n_3628);
 assign n_1979 = ~(sub_580_2_n_20 ^ n_3629);
 assign n_1981 = (sub_580_2_n_82 ^ sub_580_2_n_145);
 assign sub_580_2_n_154 = ~(sub_580_2_n_140 & (~sub_580_2_n_108 & ~sub_580_2_n_110));
 assign sub_580_2_n_153 = ~(~sub_580_2_n_33 & sub_580_2_n_149);
 assign n_1976 = ~(sub_580_2_n_18 ^ sub_580_2_n_140);
 assign sub_580_2_n_149 = ~(~sub_580_2_n_110 & sub_580_2_n_140);
 assign sub_580_2_n_145 = (~sub_580_2_n_76 | (sub_580_2_n_137 & sub_580_2_n_46));
 assign n_1980 = ~(sub_580_2_n_80 ^ sub_580_2_n_139);
 assign n_1982 = ~(sub_580_2_n_81 ^ sub_580_2_n_137);
 assign n_1983 = ~(sub_580_2_n_25 ^ n_3630);
 assign sub_580_2_n_140 = ~(~sub_580_2_n_121 & sub_580_2_n_138);
 assign sub_580_2_n_139 = ~(~sub_580_2_n_114 & sub_580_2_n_133);
 assign sub_580_2_n_138 = ~(sub_580_2_n_131 & (~sub_580_2_n_109 & ~sub_580_2_n_107));
 assign sub_580_2_n_137 = (~sub_580_2_n_103 | (sub_580_2_n_131 & sub_580_2_n_88));
 assign n_1985 = (sub_580_2_n_90 ^ sub_580_2_n_130);
 assign n_1984 = ~(sub_580_2_n_92 ^ sub_580_2_n_131);
 assign sub_580_2_n_133 = ~(~sub_580_2_n_107 & sub_580_2_n_131);
 assign sub_580_2_n_131 = ~(sub_580_2_n_128 & (~sub_580_2_n_12 & ~sub_580_2_n_111));
 assign sub_580_2_n_130 = ~(sub_580_2_n_62 & (~sub_580_2_n_60 | sub_580_2_n_127));
 assign n_1987 = (sub_580_2_n_91 ^ sub_580_2_n_37);
 assign sub_580_2_n_128 = ~(sub_580_2_n_125 & (~sub_580_2_n_95 & ~sub_580_2_n_21));
 assign sub_580_2_n_127 = ~(sub_580_2_n_106 | (~sub_580_2_n_21 & sub_580_2_n_125));
 assign n_1988 = (sub_580_2_n_23 ^ sub_580_2_n_125);
 assign sub_580_2_n_125 = ~(sub_580_2_n_123 & sub_580_2_n_8);
 assign n_1989 = (sub_580_2_n_32 ^ n_3631);
 assign sub_580_2_n_123 = ~(sub_580_2_n_79 & (sub_580_2_n_44 | (sub_580_2_n_117 & sub_580_2_n_69)));
 assign sub_580_2_n_121 = ~(sub_580_2_n_115 & (sub_580_2_n_3 & n_3632));
 assign n_1990 = ~(sub_580_2_n_117 ^ sub_580_2_n_17);
 assign sub_580_2_n_118 = ~(sub_580_2_n_113 | (~sub_580_2_n_108 & sub_580_2_n_33));
 assign sub_580_2_n_117 = ((sub_580_2_n_42 & n_572) | (n_3401 & (sub_580_2_n_42 ^ n_572)));
 assign n_1991 = (n_3401 ^ (sub_580_2_n_42 ^ n_572));
 assign sub_580_2_n_115 = ~(~sub_580_2_n_109 & sub_580_2_n_114);
 assign sub_580_2_n_114 = ~(sub_580_2_n_100 & (~sub_580_2_n_89 | sub_580_2_n_103));
 assign sub_580_2_n_113 = ~(sub_580_2_n_6 & (~sub_580_2_n_96 | sub_580_2_n_104));
 assign sub_580_2_n_111 = ~(sub_580_2_n_93 & (sub_580_2_n_105 | sub_580_2_n_95));
 assign sub_580_2_n_106 = ~sub_580_2_n_105;
 assign sub_580_2_n_110 = ~(sub_580_2_n_99 & sub_580_2_n_87);
 assign sub_580_2_n_109 = ~(sub_580_2_n_94 & sub_580_2_n_97);
 assign sub_580_2_n_108 = ~(sub_580_2_n_98 & sub_580_2_n_96);
 assign sub_580_2_n_107 = ~(sub_580_2_n_88 & sub_580_2_n_89);
 assign sub_580_2_n_105 = (~sub_580_2_n_0 & (sub_580_2_n_10 | sub_580_2_n_52));
 assign sub_580_2_n_101 = (~sub_580_2_n_5 & (sub_580_2_n_49 | sub_580_2_n_63));
 assign sub_580_2_n_100 = (~sub_580_2_n_1 & (sub_580_2_n_76 | sub_580_2_n_48));
 assign sub_580_2_n_104 = (~sub_580_2_n_16 & (sub_580_2_n_2 | sub_580_2_n_70));
 assign sub_580_2_n_103 = (~sub_580_2_n_14 & (sub_580_2_n_15 | sub_580_2_n_50));
 assign sub_580_2_n_102 = ~(sub_580_2_n_4 & (sub_580_2_n_9 | sub_580_2_n_51));
 assign sub_580_2_n_93 = ~(sub_580_2_n_61 & sub_580_2_n_65);
 assign sub_580_2_n_92 = ~(sub_580_2_n_15 & sub_580_2_n_55);
 assign sub_580_2_n_99 = ~(sub_580_2_n_47 | sub_580_2_n_53);
 assign sub_580_2_n_91 = ~(sub_580_2_n_0 | sub_580_2_n_52);
 assign sub_580_2_n_98 = ~(sub_580_2_n_66 | sub_580_2_n_70);
 assign sub_580_2_n_97 = ~(sub_580_2_n_67 | sub_580_2_n_73);
 assign sub_580_2_n_96 = ~(sub_580_2_n_57 | n_461);
 assign sub_580_2_n_95 = ~(sub_580_2_n_60 & sub_580_2_n_65);
 assign sub_580_2_n_94 = ~(sub_580_2_n_74 | sub_580_2_n_51);
 assign sub_580_2_n_90 = ~(sub_580_2_n_12 | sub_580_2_n_64);
 assign sub_580_2_n_85 = (n_623 | (n_589 | (n_410 | n_502)));
 assign n_1992 = ~(sub_580_2_n_59 & (~{in2[9]} | {in1[0]}));
 assign sub_580_2_n_83 = ~(sub_580_2_n_11 & sub_580_2_n_68);
 assign sub_580_2_n_89 = ~(sub_580_2_n_45 | sub_580_2_n_48);
 assign sub_580_2_n_82 = ~(sub_580_2_n_1 | sub_580_2_n_48);
 assign sub_580_2_n_81 = ~(sub_580_2_n_76 & sub_580_2_n_46);
 assign sub_580_2_n_88 = ~(sub_580_2_n_54 | sub_580_2_n_50);
 assign sub_580_2_n_80 = ~(sub_580_2_n_9 & sub_580_2_n_75);
 assign sub_580_2_n_87 = ~(sub_580_2_n_77 | sub_580_2_n_63);
 assign sub_580_2_n_79 = ~sub_580_2_n_78;
 assign sub_580_2_n_75 = ~sub_580_2_n_74;
 assign sub_580_2_n_72 = ~sub_580_2_n_71;
 assign sub_580_2_n_68 = ~sub_580_2_n_67;
 assign sub_580_2_n_65 = ~sub_580_2_n_64;
 assign sub_580_2_n_62 = ~sub_580_2_n_61;
 assign sub_580_2_n_78 = ~(~n_533 | n_3397);
 assign sub_580_2_n_77 = ~(~n_609 | n_3389);
 assign sub_580_2_n_76 = ~(~n_360 & n_3403);
 assign sub_580_2_n_74 = ~(~n_688 | n_3400);
 assign sub_580_2_n_73 = ~(~n_522 | n_3386);
 assign sub_580_2_n_71 = ~(~n_700 | n_3394);
 assign sub_580_2_n_70 = ~(~n_599 | n_3395);
 assign sub_580_2_n_69 = ~(sub_580_2_n_41 & n_420);
 assign sub_580_2_n_67 = ~(~n_371 | n_3390);
 assign sub_580_2_n_66 = ~(~n_481 | n_3396);
 assign sub_580_2_n_64 = ~(~n_678 | n_3388);
 assign sub_580_2_n_63 = ~(~n_451 | n_3383);
 assign sub_580_2_n_61 = ~(n_655 | sub_580_2_n_40);
 assign sub_580_2_n_60 = ~(sub_580_2_n_40 & n_655);
 assign sub_580_2_n_59 = ~({in1[0]} & ~{in2[9]});
 assign sub_580_2_n_55 = ~sub_580_2_n_54;
 assign sub_580_2_n_46 = ~sub_580_2_n_45;
 assign sub_580_2_n_43 = (n_665 | n_553);
 assign sub_580_2_n_57 = ~(~n_339 | n_3387);
 assign sub_580_2_n_56 = ~(~n_471 & n_3384);
 assign sub_580_2_n_54 = ~(~n_440 | n_3382);
 assign sub_580_2_n_53 = ~(~n_563 | n_3399);
 assign sub_580_2_n_52 = ~(~n_637 | n_3392);
 assign sub_580_2_n_51 = ~(~n_350 | n_3398);
 assign sub_580_2_n_50 = ~(~n_396 | n_3385);
 assign sub_580_2_n_49 = ~(~n_609 & n_3389);
 assign sub_580_2_n_48 = ~(~n_430 | n_3402);
 assign sub_580_2_n_47 = ~(~n_471 | n_3384);
 assign sub_580_2_n_45 = ~(~n_360 | n_3403);
 assign sub_580_2_n_44 = ~(n_420 | sub_580_2_n_41);
 assign sub_580_2_n_42 = ~n_386;
 assign sub_580_2_n_41 = ~n_3393;
 assign sub_580_2_n_40 = ~n_3391;
 assign sub_580_2_n_37 = (~sub_580_2_n_10 | (sub_580_2_n_72 & sub_580_2_n_125));
 assign sub_580_2_n_33 = ~(sub_580_2_n_101 & (~sub_580_2_n_87 | sub_580_2_n_24));
 assign sub_580_2_n_32 = ~(~sub_580_2_n_8 | sub_580_2_n_78);
 assign sub_580_2_n_31 = ~(sub_580_2_n_3 & ~sub_580_2_n_73);
 assign sub_580_2_n_30 = (sub_580_2_n_16 | sub_580_2_n_70);
 assign sub_580_2_n_29 = ~(sub_580_2_n_2 & ~sub_580_2_n_66);
 assign sub_580_2_n_28 = (sub_580_2_n_5 | sub_580_2_n_63);
 assign sub_580_2_n_27 = ~(sub_580_2_n_61 | ~sub_580_2_n_60);
 assign sub_580_2_n_26 = (sub_580_2_n_7 | sub_580_2_n_57);
 assign sub_580_2_n_25 = (sub_580_2_n_14 | sub_580_2_n_50);
 assign sub_580_2_n_24 = (sub_580_2_n_13 & (sub_580_2_n_56 | sub_580_2_n_53));
 assign sub_580_2_n_23 = ~(~sub_580_2_n_10 | sub_580_2_n_71);
 assign sub_580_2_n_22 = ~(sub_580_2_n_13 & ~sub_580_2_n_53);
 assign sub_580_2_n_21 = ~(sub_580_2_n_72 & ~sub_580_2_n_52);
 assign sub_580_2_n_20 = ~(sub_580_2_n_4 & ~sub_580_2_n_51);
 assign sub_580_2_n_19 = ~(~sub_580_2_n_49 | sub_580_2_n_77);
 assign sub_580_2_n_18 = ~(sub_580_2_n_56 & ~sub_580_2_n_47);
 assign sub_580_2_n_17 = ~(~sub_580_2_n_44 & sub_580_2_n_69);
 assign sub_580_2_n_16 = ~(n_599 | ~n_3395);
 assign sub_580_2_n_15 = ~(~n_440 & n_3382);
 assign sub_580_2_n_14 = ~(n_396 | ~n_3385);
 assign sub_580_2_n_13 = ~(~n_563 & n_3399);
 assign sub_580_2_n_12 = ~(n_678 | ~n_3388);
 assign sub_580_2_n_11 = ~(~n_371 & n_3390);
 assign sub_580_2_n_10 = ~(~n_700 & n_3394);
 assign sub_580_2_n_9 = ~(~n_688 & n_3400);
 assign sub_580_2_n_8 = ~(~n_533 & n_3397);
 assign sub_580_2_n_7 = ~(n_339 | ~n_3387);
 assign sub_580_2_n_6 = ~(sub_580_2_n_7 & ~n_461);
 assign sub_580_2_n_5 = ~(n_451 | ~n_3383);
 assign sub_580_2_n_4 = ~(~n_350 & n_3398);
 assign sub_580_2_n_3 = ~(~n_522 & n_3386);
 assign sub_580_2_n_2 = ~(~n_481 & n_3396);
 assign sub_580_2_n_1 = ~(n_430 | ~n_3402);
 assign sub_580_2_n_0 = ~(n_637 | ~n_3392);
 assign sub_599_2_n_41 = (sub_599_2_n_116 & (sub_599_2_n_39 | sub_599_2_n_106));
 assign n_2017 = ~(sub_599_2_n_99 ^ sub_599_2_n_16);
 assign n_2016 = ~(n_3152 & sub_599_2_n_171);
 assign n_2018 = (sub_599_2_n_100 ^ sub_599_2_n_41);
 assign n_2019 = ~(sub_599_2_n_35 ^ sub_599_2_n_169);
 assign n_2021 = ~(sub_599_2_n_37 ^ sub_599_2_n_170);
 assign n_2025 = (sub_599_2_n_31 ^ sub_599_2_n_168);
 assign sub_599_2_n_171 = ~(sub_599_2_n_161 | (~n_3150 | ~n_3149));
 assign sub_599_2_n_170 = ~(sub_599_2_n_15 & (sub_599_2_n_160 | sub_599_2_n_72));
 assign sub_599_2_n_169 = ~(sub_599_2_n_4 & (sub_599_2_n_39 | sub_599_2_n_63));
 assign sub_599_2_n_168 = ~(sub_599_2_n_74 | (~sub_599_2_n_60 & sub_599_2_n_159));
 assign n_2020 = (sub_599_2_n_23 ^ sub_599_2_n_39);
 assign n_2023 = (sub_599_2_n_17 ^ sub_599_2_n_26);
 assign n_2022 = (sub_599_2_n_28 ^ sub_599_2_n_160);
 assign n_2026 = ~(sub_599_2_n_21 ^ sub_599_2_n_159);
 assign n_2027 = (sub_599_2_n_30 ^ sub_599_2_n_158);
 assign n_2029 = (sub_599_2_n_27 ^ sub_599_2_n_29);
 assign sub_599_2_n_161 = ~(sub_599_2_n_36 | (sub_599_2_n_120 & (sub_599_2_n_121 & sub_599_2_n_152)));
 assign sub_599_2_n_160 = ~(sub_599_2_n_113 | (~sub_599_2_n_92 & sub_599_2_n_152));
 assign sub_599_2_n_159 = ~(sub_599_2_n_118 & (~sub_599_2_n_105 | n_3633));
 assign sub_599_2_n_158 = ~(sub_599_2_n_50 | (~sub_599_2_n_80 & sub_599_2_n_151));
 assign n_2031 = ~(sub_599_2_n_19 ^ sub_599_2_n_153);
 assign n_2024 = ~(sub_599_2_n_97 ^ sub_599_2_n_152);
 assign n_2028 = ~(sub_599_2_n_32 ^ sub_599_2_n_151);
 assign n_2030 = ~(sub_599_2_n_87 ^ sub_599_2_n_149);
 assign sub_599_2_n_153 = ~(sub_599_2_n_1 & (sub_599_2_n_145 | sub_599_2_n_81));
 assign sub_599_2_n_152 = ~(sub_599_2_n_134 & (~sub_599_2_n_123 | sub_599_2_n_145));
 assign sub_599_2_n_151 = ~n_3633;
 assign sub_599_2_n_149 = ~(sub_599_2_n_115 & (sub_599_2_n_145 | sub_599_2_n_91));
 assign n_2032 = (sub_599_2_n_33 ^ sub_599_2_n_145);
 assign n_2033 = ~(sub_599_2_n_22 ^ n_3634);
 assign sub_599_2_n_145 = ~(sub_599_2_n_139 | (~sub_599_2_n_65 | ~n_3635));
 assign n_2034 = (sub_599_2_n_20 ^ sub_599_2_n_141);
 assign n_2035 = (sub_599_2_n_24 ^ sub_599_2_n_140);
 assign sub_599_2_n_141 = ~(sub_599_2_n_112 & (~sub_599_2_n_108 | sub_599_2_n_34));
 assign sub_599_2_n_140 = ~(sub_599_2_n_3 & (~sub_599_2_n_79 | sub_599_2_n_34));
 assign sub_599_2_n_139 = ~(sub_599_2_n_34 | (~sub_599_2_n_108 | ~sub_599_2_n_95));
 assign n_2036 = (sub_599_2_n_98 ^ sub_599_2_n_34);
 assign n_2037 = ~(sub_599_2_n_101 ^ sub_599_2_n_136);
 assign sub_599_2_n_136 = ~(sub_599_2_n_13 & (sub_599_2_n_125 | sub_599_2_n_53));
 assign sub_599_2_n_135 = ~(sub_599_2_n_13 & (sub_599_2_n_53 | sub_599_2_n_125));
 assign sub_599_2_n_134 = ~(sub_599_2_n_131 | (~sub_599_2_n_84 | ~n_3636));
 assign n_2038 = (sub_599_2_n_18 ^ sub_599_2_n_125);
 assign sub_599_2_n_132 = ~(sub_599_2_n_130 & sub_599_2_n_121);
 assign sub_599_2_n_131 = ~(sub_599_2_n_129 | sub_599_2_n_119);
 assign sub_599_2_n_130 = (~sub_599_2_n_110 | (sub_599_2_n_113 & sub_599_2_n_94));
 assign sub_599_2_n_129 = ~(sub_599_2_n_109 | (sub_599_2_n_114 & sub_599_2_n_96));
 assign sub_599_2_n_127 = ~(sub_599_2_n_104 & (sub_599_2_n_116 | sub_599_2_n_93));
 assign sub_599_2_n_125 = (~n_3213 & (n_513 | sub_599_2_n_86));
 assign n_2039 = (n_513 ^ sub_599_2_n_38);
 assign sub_599_2_n_123 = ~(sub_599_2_n_122 | sub_599_2_n_119);
 assign sub_599_2_n_118 = ~sub_599_2_n_117;
 assign sub_599_2_n_122 = ~(sub_599_2_n_90 & sub_599_2_n_96);
 assign sub_599_2_n_121 = ~(sub_599_2_n_106 | sub_599_2_n_93);
 assign sub_599_2_n_120 = ~(~sub_599_2_n_94 | sub_599_2_n_92);
 assign sub_599_2_n_119 = ~(sub_599_2_n_105 & sub_599_2_n_107);
 assign sub_599_2_n_117 = ~(sub_599_2_n_0 & (sub_599_2_n_6 | sub_599_2_n_76));
 assign sub_599_2_n_115 = ~sub_599_2_n_114;
 assign sub_599_2_n_112 = ~sub_599_2_n_111;
 assign sub_599_2_n_110 = (~sub_599_2_n_2 & (sub_599_2_n_15 | sub_599_2_n_68));
 assign sub_599_2_n_109 = ~(sub_599_2_n_9 & (sub_599_2_n_75 | sub_599_2_n_71));
 assign sub_599_2_n_116 = (~sub_599_2_n_10 & (sub_599_2_n_4 | sub_599_2_n_64));
 assign sub_599_2_n_114 = ~(sub_599_2_n_11 & (sub_599_2_n_1 | sub_599_2_n_58));
 assign sub_599_2_n_113 = ~(sub_599_2_n_8 & (sub_599_2_n_70 | sub_599_2_n_52));
 assign sub_599_2_n_111 = ~(sub_599_2_n_5 & (sub_599_2_n_3 | sub_599_2_n_61));
 assign sub_599_2_n_104 = ~(sub_599_2_n_56 & sub_599_2_n_59);
 assign sub_599_2_n_101 = ~(sub_599_2_n_83 & sub_599_2_n_7);
 assign sub_599_2_n_108 = ~(sub_599_2_n_78 | sub_599_2_n_61);
 assign sub_599_2_n_107 = ~(sub_599_2_n_60 | sub_599_2_n_77);
 assign sub_599_2_n_100 = ~(sub_599_2_n_57 & sub_599_2_n_51);
 assign sub_599_2_n_106 = (sub_599_2_n_63 | sub_599_2_n_64);
 assign sub_599_2_n_99 = ~(sub_599_2_n_85 & sub_599_2_n_59);
 assign sub_599_2_n_98 = ~(sub_599_2_n_3 & sub_599_2_n_79);
 assign sub_599_2_n_105 = ~(sub_599_2_n_80 | sub_599_2_n_76);
 assign sub_599_2_n_97 = ~(sub_599_2_n_70 & sub_599_2_n_12);
 assign sub_599_2_n_91 = ~sub_599_2_n_90;
 assign n_2040 = ~(sub_599_2_n_49 & (~{in2[8]} | {in1[0]}));
 assign sub_599_2_n_87 = ~(sub_599_2_n_75 & sub_599_2_n_55);
 assign sub_599_2_n_96 = ~(sub_599_2_n_54 | sub_599_2_n_71);
 assign sub_599_2_n_95 = ~(sub_599_2_n_69 | sub_599_2_n_62);
 assign sub_599_2_n_94 = ~(sub_599_2_n_72 | sub_599_2_n_68);
 assign sub_599_2_n_93 = ~(sub_599_2_n_51 & sub_599_2_n_59);
 assign sub_599_2_n_92 = ~(~sub_599_2_n_52 & sub_599_2_n_12);
 assign sub_599_2_n_90 = ~(sub_599_2_n_81 | sub_599_2_n_58);
 assign sub_599_2_n_79 = ~sub_599_2_n_78;
 assign sub_599_2_n_74 = ~sub_599_2_n_73;
 assign sub_599_2_n_86 = ~(~n_386 | n_3425);
 assign sub_599_2_n_85 = ~(sub_599_2_n_46 & n_3409);
 assign sub_599_2_n_84 = ~(~n_522 & n_3412);
 assign sub_599_2_n_83 = ~(~n_533 & n_3420);
 assign sub_599_2_n_81 = ~(~n_440 | n_3410);
 assign sub_599_2_n_80 = ~(~n_688 | n_3424);
 assign sub_599_2_n_78 = ~(~n_700 | n_3419);
 assign sub_599_2_n_77 = ~(~n_522 | n_3412);
 assign sub_599_2_n_76 = ~(~n_350 | n_3422);
 assign sub_599_2_n_75 = ~(sub_599_2_n_43 & n_3407);
 assign sub_599_2_n_73 = ~(sub_599_2_n_44 & n_3421);
 assign sub_599_2_n_72 = ~(~n_609 | n_3415);
 assign sub_599_2_n_71 = ~(~n_430 | n_3426);
 assign sub_599_2_n_70 = ~(~n_471 & n_3408);
 assign sub_599_2_n_69 = ~(~n_655 | n_3414);
 assign sub_599_2_n_68 = ~(~n_451 | n_3411);
 assign sub_599_2_n_57 = ~sub_599_2_n_56;
 assign sub_599_2_n_55 = ~sub_599_2_n_54;
 assign sub_599_2_n_50 = ~sub_599_2_n_6;
 assign sub_599_2_n_49 = ~sub_599_2_n_48;
 assign sub_599_2_n_65 = ~(~n_678 & n_3413);
 assign sub_599_2_n_64 = ~(~n_599 | n_3418);
 assign sub_599_2_n_63 = ~(~n_481 | n_3405);
 assign sub_599_2_n_62 = ~(~n_678 | n_3413);
 assign sub_599_2_n_61 = ~(~n_637 | n_3416);
 assign sub_599_2_n_60 = ~(n_3421 | sub_599_2_n_44);
 assign sub_599_2_n_59 = (n_3409 | sub_599_2_n_46);
 assign sub_599_2_n_58 = ~(~n_396 | n_3404);
 assign sub_599_2_n_56 = ~(n_339 | sub_599_2_n_45);
 assign sub_599_2_n_54 = ~(n_3407 | sub_599_2_n_43);
 assign sub_599_2_n_53 = ~(~n_420 | n_3423);
 assign sub_599_2_n_52 = ~(~n_563 | n_3406);
 assign sub_599_2_n_51 = ~(sub_599_2_n_45 & n_339);
 assign sub_599_2_n_48 = ~({in2[8]} | ~{in1[0]});
 assign sub_599_2_n_46 = ~n_461;
 assign sub_599_2_n_45 = ~n_3417;
 assign sub_599_2_n_44 = ~n_371;
 assign sub_599_2_n_43 = ~n_360;
 assign sub_599_2_n_40 = (sub_599_2_n_120 & sub_599_2_n_152);
 assign sub_599_2_n_39 = ~(sub_599_2_n_130 | sub_599_2_n_40);
 assign sub_599_2_n_38 = (n_3213 | sub_599_2_n_86);
 assign sub_599_2_n_37 = (sub_599_2_n_2 | sub_599_2_n_68);
 assign sub_599_2_n_36 = ~(sub_599_2_n_132 & (sub_599_2_n_85 & ~sub_599_2_n_127));
 assign sub_599_2_n_35 = (sub_599_2_n_10 | sub_599_2_n_64);
 assign sub_599_2_n_34 = (sub_599_2_n_83 & ~(sub_599_2_n_135 & sub_599_2_n_7));
 assign sub_599_2_n_33 = ~(sub_599_2_n_1 & ~sub_599_2_n_81);
 assign sub_599_2_n_32 = ~(sub_599_2_n_6 & ~sub_599_2_n_80);
 assign sub_599_2_n_31 = ~(sub_599_2_n_84 & ~sub_599_2_n_77);
 assign sub_599_2_n_30 = ~(sub_599_2_n_0 & ~sub_599_2_n_76);
 assign sub_599_2_n_29 = (sub_599_2_n_75 & ~(sub_599_2_n_149 & sub_599_2_n_55));
 assign sub_599_2_n_28 = ~(sub_599_2_n_15 & ~sub_599_2_n_72);
 assign sub_599_2_n_27 = ~(sub_599_2_n_9 & ~sub_599_2_n_71);
 assign sub_599_2_n_26 = (sub_599_2_n_70 & ~(sub_599_2_n_152 & sub_599_2_n_12));
 assign sub_599_2_n_24 = ~(~sub_599_2_n_5 | sub_599_2_n_61);
 assign sub_599_2_n_23 = ~(sub_599_2_n_4 & ~sub_599_2_n_63);
 assign sub_599_2_n_22 = ~(sub_599_2_n_65 & ~sub_599_2_n_62);
 assign sub_599_2_n_21 = ~(sub_599_2_n_73 & ~sub_599_2_n_60);
 assign sub_599_2_n_20 = ~(~sub_599_2_n_14 | sub_599_2_n_69);
 assign sub_599_2_n_19 = ~(sub_599_2_n_11 & ~sub_599_2_n_58);
 assign sub_599_2_n_18 = ~(sub_599_2_n_13 & ~sub_599_2_n_53);
 assign sub_599_2_n_17 = ~(sub_599_2_n_8 & ~sub_599_2_n_52);
 assign sub_599_2_n_16 = ~(sub_599_2_n_57 & (~sub_599_2_n_51 | sub_599_2_n_41));
 assign sub_599_2_n_15 = ~(~n_609 & n_3415);
 assign sub_599_2_n_14 = ~(~n_655 & n_3414);
 assign sub_599_2_n_13 = ~(~n_420 & n_3423);
 assign sub_599_2_n_12 = ~(~n_3408 & n_471);
 assign sub_599_2_n_11 = ~(~n_396 & n_3404);
 assign sub_599_2_n_10 = ~(n_599 | ~n_3418);
 assign sub_599_2_n_9 = ~(~n_430 & n_3426);
 assign sub_599_2_n_8 = ~(~n_563 & n_3406);
 assign sub_599_2_n_7 = ~(~n_3420 & n_533);
 assign sub_599_2_n_6 = ~(~n_688 & n_3424);
 assign sub_599_2_n_5 = ~(~n_637 & n_3416);
 assign sub_599_2_n_4 = ~(~n_481 & n_3405);
 assign sub_599_2_n_3 = ~(~n_700 & n_3419);
 assign sub_599_2_n_2 = ~(n_451 | ~n_3411);
 assign sub_599_2_n_1 = ~(~n_440 & n_3410);
 assign sub_599_2_n_0 = ~(~n_350 & n_3422);
 assign n_2067 = ~(sub_618_2_n_30 ^ n_3637);
 assign n_2068 = ~(sub_618_2_n_102 ^ n_3638);
 assign n_2069 = ~(sub_618_2_n_88 ^ n_3639);
 assign n_2071 = ~(sub_618_2_n_32 ^ n_3640);
 assign n_2075 = ~(sub_618_2_n_27 ^ n_3641);
 assign n_2070 = ~(sub_618_2_n_95 ^ sub_618_2_n_174);
 assign n_2072 = ~(sub_618_2_n_93 ^ n_3652);
 assign n_2073 = ~(sub_618_2_n_31 ^ n_3642);
 assign n_2065 = ~sub_618_2_n_181;
 assign sub_618_2_n_181 = ~(sub_618_2_n_175 & sub_618_2_n_141);
 assign n_2079 = ~(sub_618_2_n_28 ^ n_3643);
 assign n_2076 = ~(sub_618_2_n_90 ^ n_3654);
 assign n_2077 = ~(sub_618_2_n_19 ^ n_3644);
 assign sub_618_2_n_175 = ~(sub_618_2_n_161 & (~sub_618_2_n_126 & ~n_3655));
 assign sub_618_2_n_174 = ~(~sub_618_2_n_33 & sub_618_2_n_170);
 assign n_2074 = ~(sub_618_2_n_89 ^ sub_618_2_n_161);
 assign sub_618_2_n_170 = ~(~sub_618_2_n_122 & sub_618_2_n_161);
 assign n_2078 = (sub_618_2_n_20 ^ n_3647);
 assign n_2080 = ~(sub_618_2_n_92 ^ n_3645);
 assign n_2081 = (sub_618_2_n_26 ^ n_3646);
 assign sub_618_2_n_161 = ~(sub_618_2_n_160 & sub_618_2_n_137);
 assign sub_618_2_n_160 = ~(sub_618_2_n_152 & (~sub_618_2_n_124 & ~sub_618_2_n_120));
 assign n_2082 = ~(sub_618_2_n_103 ^ sub_618_2_n_152);
 assign n_2083 = ~(sub_618_2_n_29 ^ n_3648);
 assign sub_618_2_n_152 = ~(sub_618_2_n_146 & (~sub_618_2_n_86 & ~sub_618_2_n_129));
 assign n_2084 = (sub_618_2_n_94 ^ n_3653);
 assign n_2085 = ~(sub_618_2_n_23 ^ n_3649);
 assign sub_618_2_n_146 = ~(sub_618_2_n_142 & (~sub_618_2_n_109 & ~sub_618_2_n_100));
 assign n_2086 = ~(sub_618_2_n_104 ^ sub_618_2_n_142);
 assign sub_618_2_n_142 = ~(~sub_618_2_n_67 & sub_618_2_n_139);
 assign sub_618_2_n_141 = ~(n_3651 | (~n_3655 & sub_618_2_n_136));
 assign n_2087 = ~(sub_618_2_n_22 ^ sub_618_2_n_138);
 assign sub_618_2_n_139 = ~(sub_618_2_n_87 & (sub_618_2_n_16 | (sub_618_2_n_134 & sub_618_2_n_58)));
 assign sub_618_2_n_138 = (sub_618_2_n_16 | (sub_618_2_n_134 & sub_618_2_n_58));
 assign sub_618_2_n_137 = ~(sub_618_2_n_131 | (~sub_618_2_n_13 | ~n_3650));
 assign sub_618_2_n_136 = ~(sub_618_2_n_132 & (~sub_618_2_n_17 & ~sub_618_2_n_127));
 assign n_2088 = (sub_618_2_n_134 ^ sub_618_2_n_91);
 assign sub_618_2_n_134 = ((sub_618_2_n_47 & n_378) | (n_926 & (sub_618_2_n_47 ^ n_378)));
 assign n_2089 = (n_926 ^ (sub_618_2_n_47 ^ n_378));
 assign sub_618_2_n_132 = ~(sub_618_2_n_33 & sub_618_2_n_123);
 assign sub_618_2_n_131 = ~(sub_618_2_n_130 | sub_618_2_n_124);
 assign sub_618_2_n_130 = ~(sub_618_2_n_114 | (sub_618_2_n_116 & sub_618_2_n_99));
 assign sub_618_2_n_129 = ~(sub_618_2_n_97 & (sub_618_2_n_118 | sub_618_2_n_100));
 assign sub_618_2_n_127 = ~((sub_618_2_n_7 | sub_618_2_n_79) & (sub_618_2_n_25 | sub_618_2_n_112));
 assign sub_618_2_n_126 = ~(~sub_618_2_n_122 & sub_618_2_n_123);
 assign sub_618_2_n_124 = ~(sub_618_2_n_111 & sub_618_2_n_108);
 assign sub_618_2_n_123 = ~(sub_618_2_n_110 | sub_618_2_n_112);
 assign sub_618_2_n_122 = ~(sub_618_2_n_113 & sub_618_2_n_101);
 assign sub_618_2_n_121 = (~sub_618_2_n_10 & (sub_618_2_n_6 | sub_618_2_n_84));
 assign sub_618_2_n_120 = ~(sub_618_2_n_107 & sub_618_2_n_99);
 assign sub_618_2_n_115 = (~sub_618_2_n_4 & (sub_618_2_n_81 | sub_618_2_n_73));
 assign sub_618_2_n_114 = ~(sub_618_2_n_18 & (sub_618_2_n_1 | sub_618_2_n_83));
 assign sub_618_2_n_118 = (~sub_618_2_n_15 & (sub_618_2_n_12 | sub_618_2_n_61));
 assign sub_618_2_n_117 = ~(sub_618_2_n_9 & (sub_618_2_n_11 | sub_618_2_n_65));
 assign sub_618_2_n_116 = ~(sub_618_2_n_5 & (sub_618_2_n_77 | sub_618_2_n_74));
 assign sub_618_2_n_113 = ~(sub_618_2_n_75 | sub_618_2_n_84);
 assign sub_618_2_n_112 = ~(sub_618_2_n_0 & sub_618_2_n_80);
 assign sub_618_2_n_104 = ~(sub_618_2_n_12 & sub_618_2_n_8);
 assign sub_618_2_n_111 = ~(sub_618_2_n_78 | sub_618_2_n_65);
 assign sub_618_2_n_110 = ~(sub_618_2_n_2 & sub_618_2_n_72);
 assign sub_618_2_n_109 = ~(sub_618_2_n_8 & sub_618_2_n_62);
 assign sub_618_2_n_103 = ~(sub_618_2_n_77 & sub_618_2_n_54);
 assign sub_618_2_n_108 = ~(sub_618_2_n_63 | sub_618_2_n_70);
 assign sub_618_2_n_107 = ~(sub_618_2_n_53 | sub_618_2_n_74);
 assign sub_618_2_n_102 = ~(sub_618_2_n_7 & sub_618_2_n_0);
 assign sub_618_2_n_97 = ~(sub_618_2_n_52 & sub_618_2_n_51);
 assign n_2090 = ~(sub_618_2_n_48 & (~{in2[7]} | {in1[0]}));
 assign sub_618_2_n_95 = ~(sub_618_2_n_69 & sub_618_2_n_2);
 assign sub_618_2_n_94 = ~(sub_618_2_n_52 | sub_618_2_n_59);
 assign sub_618_2_n_93 = ~(sub_618_2_n_81 & sub_618_2_n_50);
 assign sub_618_2_n_92 = ~(sub_618_2_n_1 & sub_618_2_n_56);
 assign sub_618_2_n_101 = ~(sub_618_2_n_49 | sub_618_2_n_73);
 assign sub_618_2_n_91 = ~(sub_618_2_n_16 | sub_618_2_n_57);
 assign sub_618_2_n_90 = ~(sub_618_2_n_82 & sub_618_2_n_64);
 assign sub_618_2_n_89 = ~(sub_618_2_n_6 & sub_618_2_n_76);
 assign sub_618_2_n_100 = ~(sub_618_2_n_60 & sub_618_2_n_51);
 assign sub_618_2_n_99 = ~(sub_618_2_n_55 | sub_618_2_n_83);
 assign sub_618_2_n_88 = ~(sub_618_2_n_3 & sub_618_2_n_72);
 assign sub_618_2_n_80 = ~sub_618_2_n_79;
 assign sub_618_2_n_76 = ~sub_618_2_n_75;
 assign sub_618_2_n_72 = ~sub_618_2_n_71;
 assign sub_618_2_n_87 = ~(sub_618_2_n_44 & n_532);
 assign sub_618_2_n_86 = ~(n_677 | sub_618_2_n_46);
 assign sub_618_2_n_84 = ~(~n_562 | n_925);
 assign sub_618_2_n_83 = ~(~n_429 | n_936);
 assign sub_618_2_n_82 = ~(sub_618_2_n_43 & n_929);
 assign sub_618_2_n_81 = ~(~n_608 & n_924);
 assign sub_618_2_n_79 = ~(~n_460 | n_914);
 assign sub_618_2_n_78 = ~(~n_687 | n_937);
 assign sub_618_2_n_77 = ~(sub_618_2_n_45 & n_915);
 assign sub_618_2_n_75 = ~(~n_470 | n_922);
 assign sub_618_2_n_74 = ~(~n_395 | n_916);
 assign sub_618_2_n_73 = ~(~n_450 | n_934);
 assign sub_618_2_n_71 = ~(~n_598 | n_923);
 assign sub_618_2_n_70 = ~(~n_521 | n_919);
 assign sub_618_2_n_69 = ~(~n_480 & n_932);
 assign sub_618_2_n_64 = ~sub_618_2_n_63;
 assign sub_618_2_n_62 = ~sub_618_2_n_61;
 assign sub_618_2_n_60 = ~sub_618_2_n_59;
 assign sub_618_2_n_58 = ~sub_618_2_n_57;
 assign sub_618_2_n_56 = ~sub_618_2_n_55;
 assign sub_618_2_n_54 = ~sub_618_2_n_53;
 assign sub_618_2_n_52 = ~sub_618_2_n_14;
 assign sub_618_2_n_50 = ~sub_618_2_n_49;
 assign sub_618_2_n_68 = ~(~n_1109 & n_2041);
 assign sub_618_2_n_67 = ~(n_532 | sub_618_2_n_44);
 assign sub_618_2_n_66 = ~(~n_1109 | n_2041);
 assign sub_618_2_n_65 = ~(~n_349 | n_920);
 assign sub_618_2_n_63 = ~(n_929 | sub_618_2_n_43);
 assign sub_618_2_n_61 = ~(~n_636 | n_935);
 assign sub_618_2_n_59 = ~(~n_654 | n_927);
 assign sub_618_2_n_57 = ~(~n_419 | n_917);
 assign sub_618_2_n_55 = ~(~n_359 | n_933);
 assign sub_618_2_n_53 = ~(n_915 | sub_618_2_n_45);
 assign sub_618_2_n_51 = ~(sub_618_2_n_46 & n_677);
 assign sub_618_2_n_49 = ~(~n_608 | n_924);
 assign sub_618_2_n_48 = ~({in1[0]} & ~{in2[7]});
 assign sub_618_2_n_47 = ~n_385;
 assign sub_618_2_n_46 = ~n_931;
 assign sub_618_2_n_45 = ~n_439;
 assign sub_618_2_n_44 = ~n_918;
 assign sub_618_2_n_43 = ~n_370;
 assign sub_618_2_n_42 = ~n_542;
 assign sub_618_2_n_33 = ~(sub_618_2_n_115 & (~sub_618_2_n_101 | sub_618_2_n_121));
 assign sub_618_2_n_32 = (sub_618_2_n_4 | sub_618_2_n_73);
 assign sub_618_2_n_31 = (sub_618_2_n_10 | sub_618_2_n_84);
 assign sub_618_2_n_30 = ~(~sub_618_2_n_17 & sub_618_2_n_80);
 assign sub_618_2_n_29 = ~(~sub_618_2_n_86 & sub_618_2_n_51);
 assign sub_618_2_n_28 = ~(sub_618_2_n_18 & ~sub_618_2_n_83);
 assign sub_618_2_n_27 = ~(sub_618_2_n_13 & ~sub_618_2_n_70);
 assign sub_618_2_n_26 = ~(~sub_618_2_n_5 | sub_618_2_n_74);
 assign sub_618_2_n_25 = (sub_618_2_n_3 & (sub_618_2_n_69 | sub_618_2_n_71));
 assign sub_618_2_n_24 = ~(~sub_618_2_n_68 | sub_618_2_n_66);
 assign sub_618_2_n_23 = ~(~sub_618_2_n_15 & sub_618_2_n_62);
 assign sub_618_2_n_22 = ~(~sub_618_2_n_67 & sub_618_2_n_87);
 assign sub_618_2_n_20 = ~(~sub_618_2_n_11 | sub_618_2_n_78);
 assign sub_618_2_n_19 = ~(sub_618_2_n_9 & ~sub_618_2_n_65);
 assign sub_618_2_n_18 = ~(~n_429 & n_936);
 assign sub_618_2_n_17 = ~(n_460 | ~n_914);
 assign sub_618_2_n_16 = ~(n_419 | ~n_917);
 assign sub_618_2_n_15 = ~(n_636 | ~n_935);
 assign sub_618_2_n_14 = ~(~n_654 & n_927);
 assign sub_618_2_n_13 = ~(~n_521 & n_919);
 assign sub_618_2_n_12 = ~(~n_699 & n_928);
 assign sub_618_2_n_11 = ~(~n_687 & n_937);
 assign sub_618_2_n_10 = ~(n_562 | ~n_925);
 assign sub_618_2_n_9 = ~(~n_349 & n_920);
 assign sub_618_2_n_8 = ~(~n_928 & n_699);
 assign sub_618_2_n_7 = ~(~n_338 & n_930);
 assign sub_618_2_n_6 = ~(~n_470 & n_922);
 assign sub_618_2_n_5 = ~(~n_395 & n_916);
 assign sub_618_2_n_4 = ~(n_450 | ~n_934);
 assign sub_618_2_n_3 = ~(~n_598 & n_923);
 assign sub_618_2_n_2 = ~(~n_932 & n_480);
 assign sub_618_2_n_1 = ~(~n_359 & n_933);
 assign sub_618_2_n_0 = ~(~n_930 & n_338);
 assign n_2122 = (sub_637_2_n_100 ^ sub_637_2_n_174);
 assign n_2119 = ~(sub_637_2_n_19 ^ n_3656);
 assign n_2117 = ~(sub_637_2_n_105 ^ n_3657);
 assign n_2120 = ~(sub_637_2_n_102 ^ sub_637_2_n_189);
 assign n_2121 = ~(sub_637_2_n_87 ^ sub_637_2_n_188);
 assign n_2123 = ~(sub_637_2_n_101 ^ n_3658);
 assign n_2127 = (sub_637_2_n_79 ^ sub_637_2_n_180);
 assign sub_637_2_n_189 = ~(sub_637_2_n_122 & (~sub_637_2_n_95 | sub_637_2_n_174));
 assign sub_637_2_n_188 = ~(sub_637_2_n_10 & (sub_637_2_n_174 | sub_637_2_n_59));
 assign n_2118 = ~(sub_637_2_n_78 ^ sub_637_2_n_175);
 assign n_2124 = ~(sub_637_2_n_85 ^ sub_637_2_n_173);
 assign n_2125 = ~(sub_637_2_n_83 ^ n_3659);
 assign n_2116 = ~(sub_637_2_n_148 | sub_637_2_n_176);
 assign sub_637_2_n_180 = ~(sub_637_2_n_60 | (~sub_637_2_n_66 & sub_637_2_n_20));
 assign n_2128 = ~(sub_637_2_n_103 ^ sub_637_2_n_20);
 assign n_2129 = ~(sub_637_2_n_98 ^ sub_637_2_n_169);
 assign n_2131 = ~(sub_637_2_n_106 ^ sub_637_2_n_168);
 assign sub_637_2_n_176 = ~(sub_637_2_n_164 | (~sub_637_2_n_128 | ~n_3664));
 assign sub_637_2_n_175 = ~(sub_637_2_n_143 & (~sub_637_2_n_128 | sub_637_2_n_164));
 assign sub_637_2_n_174 = ~(sub_637_2_n_134 | (~sub_637_2_n_22 & sub_637_2_n_163));
 assign sub_637_2_n_173 = ~(sub_637_2_n_119 & (~sub_637_2_n_112 | sub_637_2_n_164));
 assign n_2126 = ~(sub_637_2_n_80 ^ sub_637_2_n_163);
 assign sub_637_2_n_169 = ~(sub_637_2_n_56 & (n_3666 | sub_637_2_n_71));
 assign sub_637_2_n_168 = ~(sub_637_2_n_0 & (sub_637_2_n_25 | sub_637_2_n_70));
 assign n_2130 = (sub_637_2_n_82 ^ n_3666);
 assign n_2132 = (sub_637_2_n_97 ^ sub_637_2_n_25);
 assign n_2133 = ~(sub_637_2_n_104 ^ sub_637_2_n_162);
 assign sub_637_2_n_163 = ~sub_637_2_n_164;
 assign sub_637_2_n_164 = ~(sub_637_2_n_145 | (sub_637_2_n_23 & sub_637_2_n_125));
 assign sub_637_2_n_162 = ~(sub_637_2_n_7 & (sub_637_2_n_158 | sub_637_2_n_62));
 assign n_2134 = (sub_637_2_n_81 ^ sub_637_2_n_158);
 assign n_2135 = (sub_637_2_n_84 ^ sub_637_2_n_157);
 assign sub_637_2_n_158 = ~(sub_637_2_n_153 | (~sub_637_2_n_2 | ~n_3662));
 assign sub_637_2_n_157 = ~(sub_637_2_n_5 & (~sub_637_2_n_50 | sub_637_2_n_21));
 assign n_2136 = (sub_637_2_n_88 ^ sub_637_2_n_21);
 assign n_2137 = ~(sub_637_2_n_86 ^ n_3660);
 assign sub_637_2_n_153 = ~(sub_637_2_n_149 | (~sub_637_2_n_113 | ~sub_637_2_n_96));
 assign n_2138 = ~(sub_637_2_n_99 ^ sub_637_2_n_150);
 assign sub_637_2_n_150 = ~sub_637_2_n_149;
 assign sub_637_2_n_149 = ~(sub_637_2_n_57 | (sub_637_2_n_144 & sub_637_2_n_58));
 assign sub_637_2_n_148 = ~(sub_637_2_n_136 & (~n_3664 | sub_637_2_n_143));
 assign n_2139 = (sub_637_2_n_17 ^ sub_637_2_n_146);
 assign sub_637_2_n_146 = ~(sub_637_2_n_1 | (~sub_637_2_n_36 & sub_637_2_n_140));
 assign sub_637_2_n_145 = ~(sub_637_2_n_137 & (~sub_637_2_n_75 & ~sub_637_2_n_132));
 assign sub_637_2_n_144 = ~(~sub_637_2_n_1 & sub_637_2_n_141);
 assign sub_637_2_n_143 = ~(sub_637_2_n_138 | (~sub_637_2_n_6 | ~n_3663));
 assign n_2140 = ~(sub_637_2_n_140 ^ sub_637_2_n_18);
 assign sub_637_2_n_141 = ~(~sub_637_2_n_36 & sub_637_2_n_140);
 assign sub_637_2_n_140 = ((sub_618_2_n_47 & n_719) | (n_3061 & (sub_618_2_n_47 ^ n_719)));
 assign n_2141 = (n_3061 ^ (sub_618_2_n_47 ^ n_719));
 assign sub_637_2_n_138 = ~(n_3661 | sub_637_2_n_126);
 assign sub_637_2_n_137 = ~(sub_637_2_n_135 & sub_637_2_n_124);
 assign sub_637_2_n_136 = ~(sub_637_2_n_94 & (n_3153 & (sub_637_2_n_109 | sub_637_2_n_15)));
 assign sub_637_2_n_135 = (~sub_637_2_n_117 | (sub_637_2_n_118 & sub_637_2_n_92));
 assign sub_637_2_n_134 = ~n_3661;
 assign sub_637_2_n_132 = ~(sub_637_2_n_110 & (n_3665 | sub_637_2_n_111));
 assign sub_637_2_n_128 = ~(sub_637_2_n_22 | sub_637_2_n_126);
 assign sub_637_2_n_126 = ~(sub_637_2_n_95 & sub_637_2_n_114);
 assign sub_637_2_n_125 = (sub_637_2_n_115 & sub_637_2_n_92);
 assign sub_637_2_n_124 = ~(sub_637_2_n_93 | sub_637_2_n_111);
 assign sub_637_2_n_123 = ~(sub_637_2_n_76 & (sub_637_2_n_74 | sub_637_2_n_39));
 assign sub_637_2_n_122 = ~sub_637_2_n_121;
 assign sub_637_2_n_117 = (~sub_637_2_n_14 & (sub_637_2_n_0 | sub_637_2_n_67));
 assign sub_637_2_n_116 = (~sub_637_2_n_13 & (sub_637_2_n_72 | sub_637_2_n_37));
 assign sub_637_2_n_121 = ~(sub_637_2_n_12 & (sub_637_2_n_10 | sub_637_2_n_61));
 assign sub_637_2_n_119 = (~sub_637_2_n_8 & (sub_637_2_n_63 | sub_637_2_n_53));
 assign sub_637_2_n_118 = ~(sub_637_2_n_11 & (sub_637_2_n_7 | sub_637_2_n_69));
 assign sub_637_2_n_110 = ~(sub_637_2_n_60 & sub_637_2_n_38);
 assign sub_637_2_n_109 = ~(~sub_637_2_n_46 | sub_637_2_n_68);
 assign sub_637_2_n_106 = (sub_637_2_n_14 | sub_637_2_n_67);
 assign sub_637_2_n_115 = ~(sub_637_2_n_62 | sub_637_2_n_69);
 assign sub_637_2_n_105 = ~(~sub_637_2_n_15 & sub_637_2_n_46);
 assign sub_637_2_n_104 = ~(sub_637_2_n_11 & ~sub_637_2_n_69);
 assign sub_637_2_n_103 = (sub_637_2_n_60 | sub_637_2_n_66);
 assign sub_637_2_n_102 = ~(sub_637_2_n_64 & sub_637_2_n_55);
 assign sub_637_2_n_101 = (sub_637_2_n_13 | sub_637_2_n_37);
 assign sub_637_2_n_100 = ~(~sub_637_2_n_59 & sub_637_2_n_10);
 assign sub_637_2_n_99 = ~(sub_637_2_n_74 & sub_637_2_n_52);
 assign sub_637_2_n_114 = ~(sub_637_2_n_54 | sub_637_2_n_73);
 assign sub_637_2_n_113 = ~(sub_637_2_n_51 | sub_637_2_n_39);
 assign sub_637_2_n_112 = ~(sub_637_2_n_47 | sub_637_2_n_53);
 assign sub_637_2_n_98 = ~(sub_637_2_n_44 & ~sub_637_2_n_4);
 assign sub_637_2_n_111 = ~(sub_637_2_n_65 & sub_637_2_n_38);
 assign sub_637_2_n_97 = ~(sub_637_2_n_0 & ~sub_637_2_n_70);
 assign n_2142 = ~(sub_637_2_n_35 & (~{in2[6]} | {in1[0]}));
 assign sub_637_2_n_96 = ~(sub_637_2_n_49 | sub_637_2_n_42);
 assign sub_637_2_n_88 = ~(sub_637_2_n_5 & sub_637_2_n_50);
 assign sub_637_2_n_95 = ~(sub_637_2_n_59 | sub_637_2_n_61);
 assign sub_637_2_n_94 = ~(n_622 | (n_588 | (n_409 | n_501)));
 assign sub_637_2_n_87 = ~(sub_637_2_n_12 & ~sub_637_2_n_61);
 assign sub_637_2_n_93 = ~(sub_637_2_n_3 & sub_637_2_n_44);
 assign sub_637_2_n_86 = ~(sub_637_2_n_76 & ~sub_637_2_n_39);
 assign sub_637_2_n_85 = ~(sub_637_2_n_72 & sub_637_2_n_9);
 assign sub_637_2_n_84 = ~(sub_637_2_n_42 | ~sub_637_2_n_2);
 assign sub_637_2_n_83 = (sub_637_2_n_8 | sub_637_2_n_53);
 assign sub_637_2_n_82 = ~(sub_637_2_n_56 & ~sub_637_2_n_71);
 assign sub_637_2_n_81 = ~(sub_637_2_n_7 & ~sub_637_2_n_62);
 assign sub_637_2_n_80 = ~(sub_637_2_n_63 & sub_637_2_n_48);
 assign sub_637_2_n_92 = ~(sub_637_2_n_70 | sub_637_2_n_67);
 assign sub_637_2_n_79 = ~(sub_637_2_n_38 & ~sub_637_2_n_75);
 assign sub_637_2_n_78 = ~(sub_637_2_n_68 & sub_637_2_n_41);
 assign sub_637_2_n_71 = ~sub_637_2_n_3;
 assign sub_637_2_n_66 = ~sub_637_2_n_65;
 assign sub_637_2_n_76 = ~(sub_637_2_n_29 & n_3463);
 assign sub_637_2_n_75 = ~(n_521 | sub_637_2_n_30);
 assign sub_637_2_n_74 = ~(sub_637_2_n_34 & n_3466);
 assign sub_637_2_n_73 = ~(~n_460 | n_3461);
 assign sub_637_2_n_72 = ~(~n_608 & n_3453);
 assign sub_637_2_n_70 = ~(~n_359 | n_3449);
 assign sub_637_2_n_69 = ~(~n_395 | n_3457);
 assign sub_637_2_n_68 = ~(~n_1109 & n_3460);
 assign sub_637_2_n_67 = ~(~n_429 | n_2105);
 assign sub_637_2_n_65 = ~(sub_637_2_n_33 & n_370);
 assign sub_637_2_n_64 = ~(sub_637_2_n_28 & n_3450);
 assign sub_637_2_n_63 = ~(~n_470 & n_3458);
 assign sub_637_2_n_62 = ~(~n_439 | n_2108);
 assign sub_637_2_n_61 = ~(~n_598 | n_3455);
 assign sub_637_2_n_60 = ~(n_370 | sub_637_2_n_33);
 assign sub_637_2_n_59 = ~(~n_480 | n_3464);
 assign sub_637_2_n_55 = ~sub_637_2_n_54;
 assign sub_637_2_n_52 = ~sub_637_2_n_51;
 assign sub_637_2_n_50 = ~sub_637_2_n_49;
 assign sub_637_2_n_48 = ~sub_637_2_n_47;
 assign sub_637_2_n_46 = ~sub_637_2_n_45;
 assign sub_637_2_n_44 = ~sub_637_2_n_43;
 assign sub_637_2_n_41 = ~sub_637_2_n_40;
 assign sub_637_2_n_58 = ~(sub_637_2_n_32 & n_532);
 assign sub_637_2_n_57 = ~(n_532 | sub_637_2_n_32);
 assign sub_637_2_n_56 = ~(~n_687 & n_3452);
 assign sub_637_2_n_54 = ~(n_3450 | sub_637_2_n_28);
 assign sub_637_2_n_53 = ~(~n_562 | n_3456);
 assign sub_637_2_n_51 = ~(n_3466 | sub_637_2_n_34);
 assign sub_637_2_n_49 = ~(~n_654 | n_3462);
 assign sub_637_2_n_47 = ~(~n_470 | n_3458);
 assign sub_637_2_n_45 = ~(~n_542 | n_3454);
 assign sub_637_2_n_43 = ~(~n_349 | n_3469);
 assign sub_637_2_n_42 = ~(~n_677 | n_3459);
 assign sub_637_2_n_40 = ~(~n_1109 | n_3460);
 assign sub_637_2_n_39 = ~(n_3463 | sub_637_2_n_29);
 assign sub_637_2_n_38 = ~(sub_637_2_n_30 & n_521);
 assign sub_637_2_n_37 = ~(~n_450 | n_3451);
 assign sub_637_2_n_36 = ~(~n_419 | n_3060);
 assign sub_637_2_n_35 = ~({in1[0]} & ~{in2[6]});
 assign sub_637_2_n_34 = ~n_699;
 assign sub_637_2_n_33 = ~n_3467;
 assign sub_637_2_n_32 = ~n_3468;
 assign sub_637_2_n_30 = ~n_3465;
 assign sub_637_2_n_29 = ~n_636;
 assign sub_637_2_n_28 = ~n_338;
 assign sub_637_2_n_25 = ~(sub_637_2_n_118 | (~sub_637_2_n_158 & sub_637_2_n_115));
 assign sub_637_2_n_23 = ~(sub_637_2_n_158 | ~sub_637_2_n_124);
 assign sub_637_2_n_22 = ~(sub_637_2_n_112 & ~sub_637_2_n_16);
 assign sub_637_2_n_21 = ~(sub_637_2_n_123 | (sub_637_2_n_113 & sub_637_2_n_150));
 assign sub_637_2_n_20 = ~(n_3665 & (sub_637_2_n_93 | n_3666));
 assign sub_637_2_n_19 = ~(sub_637_2_n_6 & ~sub_637_2_n_73);
 assign sub_637_2_n_18 = (sub_637_2_n_1 | sub_637_2_n_36);
 assign sub_637_2_n_17 = ~(~sub_637_2_n_57 & sub_637_2_n_58);
 assign sub_637_2_n_16 = ~(sub_637_2_n_9 & ~sub_637_2_n_37);
 assign sub_637_2_n_15 = ~(n_542 | ~n_3454);
 assign sub_637_2_n_14 = ~(n_429 | ~n_2105);
 assign sub_637_2_n_13 = ~(n_450 | ~n_3451);
 assign sub_637_2_n_12 = ~(~n_598 & n_3455);
 assign sub_637_2_n_11 = ~(~n_395 & n_3457);
 assign sub_637_2_n_10 = ~(~n_480 & n_3464);
 assign sub_637_2_n_9 = ~(~n_3453 & n_608);
 assign sub_637_2_n_8 = ~(n_562 | ~n_3456);
 assign sub_637_2_n_7 = ~(~n_439 & n_2108);
 assign sub_637_2_n_6 = ~(~n_460 & n_3461);
 assign sub_637_2_n_5 = ~(~n_654 & n_3462);
 assign sub_637_2_n_4 = ~(n_349 | ~n_3469);
 assign sub_637_2_n_3 = ~(~n_3452 & n_687);
 assign sub_637_2_n_2 = ~(~n_677 & n_3459);
 assign sub_637_2_n_1 = ~(n_419 | ~n_3060);
 assign sub_637_2_n_0 = ~(~n_359 & n_3449);
 assign n_2173 = ~(n_970 ^ n_3668);
 assign n_2171 = ~(n_974 ^ n_3669);
 assign n_2170 = (n_991 ^ sub_656_2_n_27);
 assign n_2174 = ~(sub_656_2_n_90 ^ n_3670);
 assign n_2175 = ~(n_953 ^ n_3671);
 assign n_2177 = ~(n_979 ^ n_3672);
 assign n_2181 = (n_987 ^ sub_656_2_n_187);
 assign n_2172 = ~(sub_656_2_n_92 ^ n_3667);
 assign n_2176 = (n_3673 ^ sub_656_2_n_87);
 assign n_2178 = (sub_656_2_n_84 ^ n_3674);
 assign n_2179 = ~(n_1011 ^ n_3675);
 assign n_2169 = ~sub_656_2_n_188;
 assign sub_656_2_n_188 = ~(sub_656_2_n_183 & n_989);
 assign sub_656_2_n_187 = (~n_946 | (sub_656_2_n_174 & n_947));
 assign n_2182 = (sub_656_2_n_112 ^ sub_656_2_n_174);
 assign n_2183 = (n_997 ^ sub_656_2_n_173);
 assign n_2185 = ~(n_993 ^ n_3676);
 assign sub_656_2_n_183 = ~(n_1002 & (~n_976 & ~n_990));
 assign n_2180 = ~(sub_656_2_n_82 ^ n_1002);
 assign sub_656_2_n_174 = ~(n_995 & n_999);
 assign sub_656_2_n_173 = (~n_959 | (n_996 & n_998));
 assign n_2184 = ~(sub_656_2_n_93 ^ n_996);
 assign n_2186 = ~(sub_656_2_n_109 ^ n_977);
 assign n_2187 = ~(sub_656_2_n_110 ^ n_3747);
 assign sub_656_2_n_168 = ~(sub_656_2_n_164 & sub_656_2_n_98);
 assign sub_656_2_n_165 = ~(sub_656_2_n_157 & (~sub_656_2_n_130 & ~sub_656_2_n_133));
 assign sub_656_2_n_164 = ~(~sub_656_2_n_26 & sub_656_2_n_159);
 assign n_2188 = (sub_656_2_n_107 ^ sub_656_2_n_157);
 assign n_2189 = ~(sub_656_2_n_106 ^ n_3678);
 assign sub_656_2_n_159 = ~(~sub_656_2_n_133 & sub_656_2_n_157);
 assign sub_656_2_n_157 = ~(sub_656_2_n_151 & (~sub_656_2_n_80 & ~sub_656_2_n_135));
 assign n_2190 = ~(sub_656_2_n_104 ^ n_3748);
 assign n_2191 = (sub_656_2_n_103 ^ sub_656_2_n_152);
 assign sub_656_2_n_152 = (~sub_656_2_n_8 | (sub_656_2_n_148 & sub_656_2_n_2));
 assign sub_656_2_n_151 = ~(sub_656_2_n_148 & (~sub_656_2_n_17 & ~sub_656_2_n_101));
 assign n_2192 = ~(sub_656_2_n_86 ^ sub_656_2_n_148);
 assign sub_656_2_n_148 = ~(~sub_656_2_n_62 & sub_656_2_n_144);
 assign sub_656_2_n_147 = (~sub_656_2_n_145 & (sub_656_2_n_24 | n_3154));
 assign n_2193 = ~(sub_656_2_n_85 ^ sub_656_2_n_142);
 assign sub_656_2_n_145 = ~(sub_656_2_n_143 | sub_656_2_n_134);
 assign sub_656_2_n_144 = ~(sub_656_2_n_81 & (sub_656_2_n_57 | (sub_656_2_n_60 & sub_656_2_n_138)));
 assign sub_656_2_n_143 = ~(sub_656_2_n_139 | sub_656_2_n_25);
 assign sub_656_2_n_142 = (sub_656_2_n_57 | (sub_656_2_n_138 & sub_656_2_n_60));
 assign n_2194 = (sub_656_2_n_138 ^ sub_656_2_n_95);
 assign sub_656_2_n_139 = ~(sub_656_2_n_5 & (sub_656_2_n_136 | sub_656_2_n_129));
 assign sub_656_2_n_138 = ((sub_618_2_n_47 & n_571) | (n_3063 & (sub_618_2_n_47 ^ n_571)));
 assign n_2195 = (n_3063 ^ (sub_618_2_n_47 ^ n_571));
 assign sub_656_2_n_136 = (~sub_656_2_n_121 & (sub_656_2_n_127 | sub_656_2_n_116));
 assign sub_656_2_n_135 = ~(sub_656_2_n_114 & (sub_656_2_n_125 | sub_656_2_n_101));
 assign sub_656_2_n_134 = ~(sub_656_2_n_120 & (~n_3154 & ~sub_656_2_n_18));
 assign sub_656_2_n_133 = ~(sub_656_2_n_99 & sub_656_2_n_119);
 assign sub_656_2_n_132 = ~(sub_656_2_n_118 | sub_656_2_n_116);
 assign sub_656_2_n_130 = ~(sub_656_2_n_98 & sub_656_2_n_102);
 assign sub_656_2_n_129 = ~(sub_656_2_n_100 & sub_656_2_n_117);
 assign sub_656_2_n_128 = (~sub_656_2_n_3 & (sub_656_2_n_42 | sub_656_2_n_73));
 assign sub_656_2_n_127 = (~sub_656_2_n_16 & (sub_656_2_n_68 | sub_656_2_n_58));
 assign sub_656_2_n_122 = (~sub_656_2_n_4 & (sub_656_2_n_72 | sub_656_2_n_79));
 assign sub_656_2_n_121 = ~(sub_656_2_n_10 & (sub_656_2_n_11 | sub_656_2_n_59));
 assign sub_656_2_n_126 = (~sub_656_2_n_6 & (sub_656_2_n_55 | sub_656_2_n_44));
 assign sub_656_2_n_125 = (~sub_656_2_n_15 & (sub_656_2_n_8 | sub_656_2_n_46));
 assign sub_656_2_n_124 = ~(sub_656_2_n_0 & (~sub_656_2_n_13 | sub_656_2_n_52));
 assign sub_656_2_n_123 = (~sub_656_2_n_1 & (sub_656_2_n_56 | sub_656_2_n_45));
 assign sub_656_2_n_115 = ~(sub_656_2_n_7 & sub_656_2_n_41);
 assign sub_656_2_n_114 = ~(sub_656_2_n_77 & sub_656_2_n_76);
 assign sub_656_2_n_113 = ~(sub_656_2_n_63 | n_552);
 assign sub_656_2_n_120 = ~(~sub_656_2_n_13 | sub_656_2_n_66);
 assign sub_656_2_n_112 = (n_946 & n_947);
 assign sub_656_2_n_111 = ~(sub_656_2_n_6 | sub_656_2_n_44);
 assign sub_656_2_n_110 = (sub_656_2_n_3 | sub_656_2_n_73);
 assign sub_656_2_n_109 = ~(n_983 & n_982);
 assign sub_656_2_n_108 = ~(sub_656_2_n_12 | sub_656_2_n_67);
 assign sub_656_2_n_119 = ~(sub_656_2_n_74 | sub_656_2_n_79);
 assign sub_656_2_n_107 = (sub_656_2_n_42 & sub_656_2_n_51);
 assign sub_656_2_n_106 = ~(~sub_656_2_n_80 & sub_656_2_n_76);
 assign sub_656_2_n_105 = ~(sub_656_2_n_10 & ~sub_656_2_n_59);
 assign sub_656_2_n_104 = ~(sub_656_2_n_78 & sub_656_2_n_39);
 assign sub_656_2_n_103 = ~(sub_656_2_n_15 | sub_656_2_n_46);
 assign sub_656_2_n_118 = ~(~sub_656_2_n_58 & sub_656_2_n_9);
 assign sub_656_2_n_117 = ~(sub_656_2_n_53 | sub_656_2_n_40);
 assign sub_656_2_n_116 = (sub_656_2_n_65 | sub_656_2_n_59);
 assign n_2196 = ~(sub_656_2_n_64 & (~{in2[5]} | {in1[0]}));
 assign sub_656_2_n_102 = ~(sub_656_2_n_48 | sub_656_2_n_67);
 assign sub_656_2_n_95 = ~(~sub_656_2_n_60 | sub_656_2_n_57);
 assign sub_656_2_n_94 = ~(sub_656_2_n_0 & sub_656_2_n_13);
 assign sub_656_2_n_93 = ~(n_959 & n_998);
 assign sub_656_2_n_92 = ~(~n_966 & n_1015);
 assign sub_656_2_n_101 = ~(sub_656_2_n_39 & sub_656_2_n_76);
 assign sub_656_2_n_91 = ~(sub_656_2_n_5 & sub_656_2_n_41);
 assign sub_656_2_n_90 = ~(n_940 & n_942);
 assign sub_656_2_n_89 = (sub_656_2_n_1 | sub_656_2_n_45);
 assign sub_656_2_n_88 = (sub_656_2_n_4 | sub_656_2_n_79);
 assign sub_656_2_n_87 = ~(~n_944 | n_943);
 assign sub_656_2_n_86 = ~(sub_656_2_n_8 & sub_656_2_n_2);
 assign sub_656_2_n_100 = ~(sub_656_2_n_71 | sub_656_2_n_45);
 assign sub_656_2_n_85 = ~(~sub_656_2_n_62 & sub_656_2_n_81);
 assign sub_656_2_n_84 = ~(n_1005 | ~n_962);
 assign sub_656_2_n_83 = (sub_656_2_n_16 | sub_656_2_n_58);
 assign sub_656_2_n_99 = ~(sub_656_2_n_50 | sub_656_2_n_73);
 assign sub_656_2_n_82 = ~(n_1013 & n_980);
 assign sub_656_2_n_98 = ~(sub_656_2_n_69 | sub_656_2_n_44);
 assign sub_656_2_n_78 = ~sub_656_2_n_77;
 assign sub_656_2_n_75 = ~sub_656_2_n_74;
 assign sub_656_2_n_70 = ~sub_656_2_n_69;
 assign sub_656_2_n_81 = ~(sub_656_2_n_37 & n_532);
 assign sub_656_2_n_80 = ~(n_677 | sub_656_2_n_32);
 assign sub_656_2_n_79 = ~(~n_429 | n_3476);
 assign sub_656_2_n_77 = ~(n_654 | sub_656_2_n_34);
 assign sub_656_2_n_76 = ~(sub_656_2_n_32 & n_677);
 assign sub_656_2_n_74 = ~(~n_359 | n_3479);
 assign sub_656_2_n_73 = ~(~n_395 | n_2160);
 assign sub_656_2_n_72 = ~(~n_359 & n_3479);
 assign sub_656_2_n_71 = ~(~n_480 | n_3472);
 assign sub_656_2_n_69 = ~(~n_687 | n_3475);
 assign sub_656_2_n_68 = ~(~n_470 & n_3487);
 assign sub_656_2_n_67 = ~(~n_521 | n_3489);
 assign sub_656_2_n_66 = ~(n_3483 | sub_656_2_n_38);
 assign sub_656_2_n_65 = ~(~n_608 | n_3478);
 assign sub_656_2_n_64 = ~({in1[0]} & ~{in2[5]});
 assign sub_656_2_n_54 = ~sub_656_2_n_53;
 assign sub_656_2_n_51 = ~sub_656_2_n_50;
 assign sub_656_2_n_49 = ~sub_656_2_n_48;
 assign sub_656_2_n_47 = ~sub_656_2_n_14;
 assign sub_656_2_n_43 = ~sub_656_2_n_7;
 assign sub_656_2_n_41 = ~sub_656_2_n_40;
 assign sub_656_2_n_63 = ~(sub_656_2_n_33 & n_3470);
 assign sub_656_2_n_62 = ~(n_532 | sub_656_2_n_37);
 assign sub_656_2_n_61 = ~(n_3470 | sub_656_2_n_33);
 assign sub_656_2_n_60 = ~(sub_656_2_n_35 & n_419);
 assign sub_656_2_n_59 = ~(~n_450 | n_3474);
 assign sub_656_2_n_58 = ~(~n_562 | n_3480);
 assign sub_656_2_n_57 = ~(n_419 | sub_656_2_n_35);
 assign sub_656_2_n_56 = ~(~n_480 & n_3472);
 assign sub_656_2_n_55 = ~(~n_687 & n_3475);
 assign sub_656_2_n_53 = ~(~n_338 | n_3477);
 assign sub_656_2_n_52 = ~(sub_656_2_n_38 & n_3483);
 assign sub_656_2_n_50 = ~(~n_439 | n_3481);
 assign sub_656_2_n_48 = ~(~n_370 | n_3491);
 assign sub_656_2_n_46 = ~(~n_636 | n_3488);
 assign sub_656_2_n_45 = ~(~n_598 | n_3486);
 assign sub_656_2_n_44 = ~(~n_349 | n_3473);
 assign sub_656_2_n_42 = ~(~n_439 & n_3481);
 assign sub_656_2_n_40 = ~(~n_460 | n_3471);
 assign sub_656_2_n_39 = ~(sub_656_2_n_34 & n_654);
 assign sub_656_2_n_38 = ~n_1109;
 assign sub_656_2_n_37 = ~n_2166;
 assign sub_656_2_n_35 = ~n_3062;
 assign sub_656_2_n_34 = ~n_3485;
 assign sub_656_2_n_33 = ~n_664;
 assign sub_656_2_n_32 = ~n_3484;
 assign sub_656_2_n_29 = ~(sub_656_2_n_132 & ~sub_656_2_n_129);
 assign sub_656_2_n_27 = (n_965 | (n_3667 & n_973));
 assign sub_656_2_n_26 = ~(sub_656_2_n_122 & (~sub_656_2_n_119 | sub_656_2_n_128));
 assign sub_656_2_n_25 = ~(sub_656_2_n_115 & (~sub_656_2_n_117 | sub_656_2_n_123));
 assign sub_656_2_n_24 = ~(sub_656_2_n_113 | (~sub_656_2_n_18 & sub_656_2_n_124));
 assign sub_656_2_n_23 = ~(sub_656_2_n_20 & (~sub_656_2_n_102 | sub_656_2_n_126));
 assign sub_656_2_n_20 = ~(sub_656_2_n_14 & ~sub_656_2_n_67);
 assign sub_656_2_n_19 = ~(~sub_656_2_n_63 | sub_656_2_n_61);
 assign sub_656_2_n_18 = (n_552 | sub_656_2_n_61);
 assign sub_656_2_n_17 = ~(sub_656_2_n_2 & ~sub_656_2_n_46);
 assign sub_656_2_n_16 = ~(n_562 | ~n_3480);
 assign sub_656_2_n_15 = ~(n_636 | ~n_3488);
 assign sub_656_2_n_14 = ~(n_370 | ~n_3491);
 assign sub_656_2_n_13 = ~(~n_3482 & n_542);
 assign sub_656_2_n_12 = ~(n_521 | ~n_3489);
 assign sub_656_2_n_11 = ~(~n_608 & n_3478);
 assign sub_656_2_n_10 = ~(~n_450 & n_3474);
 assign sub_656_2_n_9 = ~(~n_3487 & n_470);
 assign sub_656_2_n_8 = ~(~n_699 & n_3490);
 assign sub_656_2_n_7 = ~(n_338 | ~n_3477);
 assign sub_656_2_n_6 = ~(n_349 | ~n_3473);
 assign sub_656_2_n_5 = ~(~n_460 & n_3471);
 assign sub_656_2_n_4 = ~(n_429 | ~n_3476);
 assign sub_656_2_n_3 = ~(n_395 | ~n_2160);
 assign sub_656_2_n_2 = ~(~n_3490 & n_699);
 assign sub_656_2_n_1 = ~(n_598 | ~n_3486);
 assign sub_656_2_n_0 = ~(~n_542 & n_3482);
 assign sub_675_2_n_19 = (n_3685 & ~(n_3181 & sub_675_2_n_119));
 assign n_2225 = ~(sub_675_2_n_73 ^ sub_675_2_n_207);
 assign n_2229 = ~(sub_675_2_n_80 ^ sub_675_2_n_15);
 assign sub_675_2_n_207 = ~(sub_675_2_n_67 & (sub_675_2_n_19 | sub_675_2_n_48));
 assign n_2226 = ~(sub_675_2_n_83 ^ sub_675_2_n_19);
 assign n_2227 = ~(sub_675_2_n_82 ^ sub_675_2_n_198);
 assign n_2230 = ~(sub_675_2_n_79 ^ sub_675_2_n_197);
 assign n_2231 = ~(sub_675_2_n_102 ^ sub_675_2_n_196);
 assign n_2233 = ~(sub_675_2_n_75 ^ n_3679);
 assign n_2224 = ~(sub_675_2_n_144 | sub_675_2_n_199);
 assign n_2237 = ~(sub_675_2_n_14 ^ sub_675_2_n_188);
 assign sub_675_2_n_199 = ~(sub_675_2_n_128 | sub_675_2_n_189);
 assign sub_675_2_n_198 = (~sub_675_2_n_60 | (n_3181 & sub_675_2_n_54));
 assign sub_675_2_n_197 = ~(sub_675_2_n_127 | (sub_675_2_n_181 & sub_675_2_n_91));
 assign sub_675_2_n_196 = (~sub_675_2_n_0 | (sub_675_2_n_181 & sub_675_2_n_3));
 assign n_2235 = ~(sub_675_2_n_84 ^ sub_675_2_n_184);
 assign n_2228 = ~(sub_675_2_n_81 ^ n_3181);
 assign n_2232 = ~(sub_675_2_n_77 ^ sub_675_2_n_181);
 assign n_2234 = ~(sub_675_2_n_74 ^ n_3680);
 assign sub_675_2_n_189 = ~(~sub_675_2_n_94 & n_3181);
 assign sub_675_2_n_188 = ~(sub_675_2_n_1 & (sub_675_2_n_16 | sub_675_2_n_42));
 assign n_2238 = (sub_675_2_n_108 ^ sub_675_2_n_16);
 assign n_2239 = ~(sub_675_2_n_106 ^ sub_675_2_n_175);
 assign n_2241 = ~(sub_675_2_n_107 ^ sub_675_2_n_174);
 assign sub_675_2_n_184 = ~(sub_675_2_n_40 & (sub_675_2_n_170 | sub_675_2_n_36));
 assign sub_675_2_n_181 = ~(~sub_675_2_n_17 & sub_675_2_n_176);
 assign n_2236 = ~(sub_675_2_n_104 ^ sub_675_2_n_170);
 assign sub_675_2_n_176 = ~(~sub_675_2_n_131 & sub_675_2_n_169);
 assign sub_675_2_n_175 = (~sub_675_2_n_5 | (n_3681 & sub_675_2_n_65));
 assign sub_675_2_n_174 = ~(sub_675_2_n_7 & (sub_675_2_n_166 | sub_675_2_n_63));
 assign n_2240 = ~(sub_675_2_n_105 ^ n_3681);
 assign n_2242 = (sub_675_2_n_103 ^ sub_675_2_n_166);
 assign n_2243 = ~(sub_675_2_n_109 ^ sub_675_2_n_165);
 assign sub_675_2_n_170 = ~sub_675_2_n_169;
 assign sub_675_2_n_169 = ~(~sub_675_2_n_146 & sub_675_2_n_168);
 assign sub_675_2_n_168 = ~(n_3177 & (~sub_675_2_n_129 & ~sub_675_2_n_132));
 assign sub_675_2_n_166 = ~(sub_675_2_n_130 | (n_3177 & sub_675_2_n_118));
 assign sub_675_2_n_165 = (~sub_675_2_n_10 | (n_3177 & sub_675_2_n_35));
 assign n_2244 = ~(n_3177 ^ sub_675_2_n_98);
 assign n_2245 = (sub_675_2_n_76 ^ sub_675_2_n_159);
 assign sub_675_2_n_159 = ~(sub_675_2_n_61 | (sub_675_2_n_156 & sub_675_2_n_30));
 assign n_2246 = ~(sub_675_2_n_101 ^ sub_675_2_n_156);
 assign n_2247 = ~(sub_675_2_n_78 ^ sub_675_2_n_155);
 assign sub_675_2_n_156 = ~(sub_675_2_n_123 & (sub_675_2_n_151 | sub_675_2_n_95));
 assign sub_675_2_n_155 = ~(sub_675_2_n_9 & (sub_675_2_n_151 | sub_675_2_n_57));
 assign sub_675_2_n_154 = ~(sub_675_2_n_152 & (~sub_675_2_n_117 & ~sub_675_2_n_95));
 assign n_2248 = ~((sub_675_2_n_151 & ~sub_675_2_n_100) | (sub_675_2_n_152 & sub_675_2_n_100));
 assign sub_675_2_n_151 = ~sub_675_2_n_152;
 assign sub_675_2_n_152 = ~(sub_675_2_n_149 & sub_675_2_n_50);
 assign n_2249 = (sub_675_2_n_99 ^ sub_675_2_n_147);
 assign sub_675_2_n_149 = ~(n_3214 & (sub_675_2_n_41 | (sub_675_2_n_143 & sub_675_2_n_49)));
 assign sub_675_2_n_148 = ~(sub_675_2_n_141 & (~sub_675_2_n_69 & ~sub_675_2_n_137));
 assign sub_675_2_n_147 = ~(sub_675_2_n_41 | (sub_675_2_n_143 & sub_675_2_n_49));
 assign sub_675_2_n_146 = ~(sub_675_2_n_4 & (n_3682 & (sub_675_2_n_139 | sub_675_2_n_132)));
 assign n_2250 = ~(sub_675_2_n_143 ^ sub_675_2_n_85);
 assign sub_675_2_n_144 = ~(sub_675_2_n_140 | sub_675_2_n_89);
 assign sub_675_2_n_143 = ((sub_694_2_n_13 & n_380) | (n_3064 & (sub_694_2_n_13 ^ n_380)));
 assign n_2251 = (n_3064 ^ (sub_694_2_n_13 ^ n_380));
 assign sub_675_2_n_141 = ~(sub_675_2_n_17 & sub_675_2_n_133);
 assign sub_675_2_n_140 = ~(sub_675_2_n_134 | (~sub_675_2_n_87 | ~sub_675_2_n_51));
 assign sub_675_2_n_139 = ~(sub_675_2_n_121 | (sub_675_2_n_115 & sub_675_2_n_130));
 assign sub_675_2_n_138 = ~(sub_675_2_n_110 & (sub_675_2_n_123 | sub_675_2_n_117));
 assign sub_675_2_n_137 = ~(sub_675_2_n_111 & (sub_675_2_n_126 | sub_675_2_n_97));
 assign sub_675_2_n_135 = ~(~sub_675_2_n_131 & sub_675_2_n_133);
 assign sub_675_2_n_134 = ~(n_3685 | sub_675_2_n_94);
 assign sub_675_2_n_128 = ~(~sub_675_2_n_89 & sub_675_2_n_119);
 assign sub_675_2_n_133 = ~(sub_675_2_n_90 | sub_675_2_n_97);
 assign sub_675_2_n_132 = ~(sub_675_2_n_92 & sub_675_2_n_96);
 assign sub_675_2_n_131 = ~(sub_675_2_n_116 & sub_675_2_n_93);
 assign sub_675_2_n_130 = ~(sub_675_2_n_70 & (sub_675_2_n_10 | sub_675_2_n_32));
 assign sub_675_2_n_129 = ~(sub_675_2_n_118 & sub_675_2_n_115);
 assign sub_675_2_n_127 = ~sub_675_2_n_126;
 assign sub_675_2_n_121 = ~(sub_675_2_n_2 & (sub_675_2_n_7 | sub_675_2_n_56));
 assign sub_675_2_n_126 = (~sub_675_2_n_8 & (sub_675_2_n_0 | sub_675_2_n_45));
 assign sub_675_2_n_125 = ~(sub_675_2_n_13 & (sub_675_2_n_5 | sub_675_2_n_37));
 assign sub_675_2_n_123 = (~sub_675_2_n_11 & (sub_675_2_n_9 | sub_675_2_n_31));
 assign sub_675_2_n_111 = ~(sub_675_2_n_55 & sub_675_2_n_58);
 assign sub_675_2_n_110 = ~(sub_675_2_n_61 & sub_675_2_n_62);
 assign sub_675_2_n_109 = ~(sub_675_2_n_70 & ~sub_675_2_n_32);
 assign sub_675_2_n_108 = ~(sub_675_2_n_1 & ~sub_675_2_n_42);
 assign sub_675_2_n_107 = ~(sub_675_2_n_2 & ~sub_675_2_n_56);
 assign sub_675_2_n_106 = ~(sub_675_2_n_13 & ~sub_675_2_n_37);
 assign sub_675_2_n_119 = ~(sub_675_2_n_53 | sub_675_2_n_59);
 assign sub_675_2_n_118 = ~(sub_675_2_n_34 | sub_675_2_n_32);
 assign sub_675_2_n_105 = ~(sub_675_2_n_5 & sub_675_2_n_65);
 assign sub_675_2_n_104 = ~(~sub_675_2_n_40 | sub_675_2_n_36);
 assign sub_675_2_n_103 = ~(sub_675_2_n_7 & ~sub_675_2_n_63);
 assign sub_675_2_n_117 = ~(sub_675_2_n_30 & sub_675_2_n_62);
 assign sub_675_2_n_102 = (sub_675_2_n_8 | sub_675_2_n_45);
 assign sub_675_2_n_101 = ~(sub_675_2_n_30 & ~sub_675_2_n_61);
 assign sub_675_2_n_100 = ~(~sub_675_2_n_9 | sub_675_2_n_57);
 assign sub_675_2_n_99 = ~(sub_675_2_n_50 & n_3214);
 assign sub_675_2_n_116 = ~(sub_675_2_n_36 | sub_675_2_n_33);
 assign sub_675_2_n_98 = ~(sub_675_2_n_10 & sub_675_2_n_35);
 assign sub_675_2_n_115 = ~(sub_675_2_n_63 | sub_675_2_n_56);
 assign sub_675_2_n_91 = ~sub_675_2_n_90;
 assign sub_675_2_n_87 = ~(~sub_675_2_n_67 & sub_675_2_n_66);
 assign n_2252 = ~(sub_675_2_n_29 & (~{in2[4]} | {in1[0]}));
 assign sub_675_2_n_85 = ~(sub_675_2_n_49 & ~sub_675_2_n_41);
 assign sub_675_2_n_97 = ~(sub_675_2_n_43 & sub_675_2_n_58);
 assign sub_675_2_n_96 = ~(sub_675_2_n_42 | sub_675_2_n_47);
 assign sub_675_2_n_84 = (sub_675_2_n_6 | sub_675_2_n_33);
 assign sub_675_2_n_83 = ~(~sub_675_2_n_67 | sub_675_2_n_48);
 assign sub_675_2_n_95 = (sub_675_2_n_57 | sub_675_2_n_31);
 assign sub_675_2_n_82 = (sub_675_2_n_72 | sub_675_2_n_59);
 assign sub_675_2_n_81 = ~(sub_675_2_n_60 & sub_675_2_n_54);
 assign sub_675_2_n_94 = ~(~sub_675_2_n_48 & sub_675_2_n_66);
 assign sub_675_2_n_80 = ~(~sub_675_2_n_69 & sub_675_2_n_58);
 assign sub_675_2_n_93 = ~(sub_675_2_n_38 | sub_675_2_n_46);
 assign sub_675_2_n_79 = ~(sub_675_2_n_55 | sub_675_2_n_44);
 assign sub_675_2_n_92 = ~(sub_675_2_n_64 | sub_675_2_n_37);
 assign sub_675_2_n_78 = (sub_675_2_n_11 | sub_675_2_n_31);
 assign sub_675_2_n_77 = ~(sub_675_2_n_0 & sub_675_2_n_3);
 assign sub_675_2_n_76 = ~(sub_675_2_n_62 & ~sub_675_2_n_52);
 assign sub_675_2_n_75 = ~(sub_675_2_n_12 & ~sub_675_2_n_46);
 assign sub_675_2_n_90 = ~(~sub_675_2_n_45 & sub_675_2_n_3);
 assign sub_675_2_n_74 = ~(sub_675_2_n_68 & sub_675_2_n_39);
 assign sub_675_2_n_73 = ~(sub_675_2_n_51 & sub_675_2_n_66);
 assign sub_675_2_n_89 = (n_621 | (n_587 | (n_408 | n_500)));
 assign sub_675_2_n_65 = ~sub_675_2_n_64;
 assign sub_675_2_n_54 = ~sub_675_2_n_53;
 assign sub_675_2_n_72 = ~(n_541 | ~n_3505);
 assign sub_675_2_n_70 = ~(sub_675_2_n_26 & n_3514);
 assign sub_675_2_n_69 = ~(n_459 | sub_675_2_n_22);
 assign sub_675_2_n_68 = ~(~n_607 & n_3503);
 assign sub_675_2_n_67 = ~(~n_663 & n_3504);
 assign sub_675_2_n_66 = ~(n_551 & ~n_3492);
 assign sub_675_2_n_64 = ~(~n_686 | n_3498);
 assign sub_675_2_n_63 = ~(~n_358 | n_3502);
 assign sub_675_2_n_62 = ~(sub_675_2_n_25 & n_676);
 assign sub_675_2_n_61 = ~(n_653 | sub_675_2_n_21);
 assign sub_675_2_n_60 = ~(~n_1108 & n_3493);
 assign sub_675_2_n_59 = ~(~n_541 | n_3505);
 assign sub_675_2_n_58 = ~(sub_675_2_n_22 & n_459);
 assign sub_675_2_n_57 = ~(~n_698 | n_3067);
 assign sub_675_2_n_56 = ~(~n_428 | n_3501);
 assign sub_675_2_n_55 = ~(n_337 | sub_675_2_n_28);
 assign sub_675_2_n_53 = ~(~n_1108 | n_3493);
 assign sub_675_2_n_44 = ~sub_675_2_n_43;
 assign sub_675_2_n_39 = ~sub_675_2_n_38;
 assign sub_675_2_n_35 = ~sub_675_2_n_34;
 assign sub_675_2_n_52 = ~(n_676 | sub_675_2_n_25);
 assign sub_675_2_n_51 = ~(~n_551 & n_3492);
 assign sub_675_2_n_50 = ~(~n_531 & n_3513);
 assign sub_675_2_n_49 = ~(sub_675_2_n_24 & n_418);
 assign sub_675_2_n_48 = ~(~n_663 | n_3504);
 assign sub_675_2_n_47 = ~(~n_520 | n_3512);
 assign sub_675_2_n_46 = ~(~n_449 | n_3500);
 assign sub_675_2_n_45 = ~(~n_597 | n_3494);
 assign sub_675_2_n_43 = ~(sub_675_2_n_28 & n_337);
 assign sub_675_2_n_42 = ~(~n_369 | n_3495);
 assign sub_675_2_n_41 = ~(n_418 | sub_675_2_n_24);
 assign sub_675_2_n_40 = ~(~n_469 & n_3510);
 assign sub_675_2_n_38 = ~(~n_607 | n_3503);
 assign sub_675_2_n_37 = ~(~n_348 | n_3497);
 assign sub_675_2_n_36 = ~(~n_469 | n_3510);
 assign sub_675_2_n_34 = ~(~n_438 | n_3066);
 assign sub_675_2_n_33 = ~(~n_561 | n_3508);
 assign sub_675_2_n_32 = ~(n_3514 | sub_675_2_n_26);
 assign sub_675_2_n_31 = ~(~n_635 | n_3511);
 assign sub_675_2_n_30 = ~(sub_675_2_n_21 & n_653);
 assign sub_675_2_n_29 = ~({in1[0]} & ~{in2[4]});
 assign sub_675_2_n_28 = ~n_3507;
 assign sub_675_2_n_26 = ~n_394;
 assign sub_675_2_n_25 = ~n_3506;
 assign sub_675_2_n_24 = ~n_3065;
 assign sub_675_2_n_22 = ~n_3499;
 assign sub_675_2_n_21 = ~n_3509;
 assign sub_675_2_n_17 = ~(n_3683 & (~sub_675_2_n_93 | n_3684));
 assign sub_675_2_n_16 = ~(sub_675_2_n_125 | (sub_675_2_n_92 & n_3681));
 assign sub_675_2_n_15 = ~(~sub_675_2_n_55 & (sub_675_2_n_197 | sub_675_2_n_44));
 assign sub_675_2_n_14 = ~(sub_675_2_n_4 & ~sub_675_2_n_47);
 assign sub_675_2_n_13 = ~(~n_348 & n_3497);
 assign sub_675_2_n_12 = ~(~n_449 & n_3500);
 assign sub_675_2_n_11 = ~(n_635 | ~n_3511);
 assign sub_675_2_n_10 = ~(~n_438 & n_3066);
 assign sub_675_2_n_9 = ~(~n_698 & n_3067);
 assign sub_675_2_n_8 = ~(n_597 | ~n_3494);
 assign sub_675_2_n_7 = ~(~n_358 & n_3502);
 assign sub_675_2_n_6 = ~(n_561 | ~n_3508);
 assign sub_675_2_n_5 = ~(~n_686 & n_3498);
 assign sub_675_2_n_4 = ~(~n_520 & n_3512);
 assign sub_675_2_n_3 = ~(~n_3496 & n_479);
 assign sub_675_2_n_2 = ~(~n_428 & n_3501);
 assign sub_675_2_n_1 = ~(~n_369 & n_3495);
 assign sub_675_2_n_0 = ~(~n_479 & n_3496);
 assign sub_694_2_n_7 = ~(sub_694_2_n_110 | (~sub_694_2_n_176 & sub_694_2_n_102));
 assign n_2283 = (sub_694_2_n_75 ^ sub_694_2_n_196);
 assign n_2287 = (sub_694_2_n_70 ^ sub_694_2_n_192);
 assign sub_694_2_n_196 = ~(sub_694_2_n_28 & (sub_694_2_n_7 | sub_694_2_n_26));
 assign n_2282 = (sub_694_2_n_64 ^ sub_694_2_n_188);
 assign n_2284 = (sub_694_2_n_98 ^ sub_694_2_n_7);
 assign n_2285 = (sub_694_2_n_87 ^ sub_694_2_n_187);
 assign sub_694_2_n_192 = ~(sub_694_2_n_53 & (sub_694_2_n_183 | sub_694_2_n_30));
 assign n_2291 = ~(sub_694_2_n_86 ^ sub_694_2_n_184);
 assign n_2288 = ~(sub_694_2_n_68 ^ sub_694_2_n_183);
 assign n_2289 = ~(sub_694_2_n_67 ^ sub_694_2_n_182);
 assign sub_694_2_n_188 = ~(sub_694_2_n_129 & (sub_694_2_n_176 | sub_694_2_n_122));
 assign sub_694_2_n_187 = ~(sub_694_2_n_43 & (sub_694_2_n_176 | sub_694_2_n_21));
 assign n_2295 = ~(sub_694_2_n_92 ^ sub_694_2_n_175);
 assign n_2286 = (sub_694_2_n_71 ^ sub_694_2_n_176);
 assign sub_694_2_n_184 = ~(sub_694_2_n_1 & (sub_694_2_n_171 | sub_694_2_n_40));
 assign sub_694_2_n_183 = ~(sub_694_2_n_113 | (sub_694_2_n_168 & sub_694_2_n_103));
 assign sub_694_2_n_182 = (~sub_694_2_n_24 | (sub_694_2_n_168 & sub_694_2_n_4));
 assign n_2292 = ~(sub_694_2_n_72 ^ sub_694_2_n_171);
 assign n_2293 = ~(sub_694_2_n_97 ^ sub_694_2_n_170);
 assign n_2290 = ~(sub_694_2_n_65 ^ sub_694_2_n_168);
 assign sub_694_2_n_176 = (sub_694_2_n_169 & sub_694_2_n_136);
 assign sub_694_2_n_175 = ~(sub_694_2_n_15 & (sub_694_2_n_166 | sub_694_2_n_23));
 assign n_2296 = ~(sub_694_2_n_95 ^ sub_694_2_n_166);
 assign n_2297 = ~(sub_694_2_n_99 ^ sub_694_2_n_165);
 assign n_2299 = ~(sub_694_2_n_89 ^ sub_694_2_n_164);
 assign sub_694_2_n_171 = ~(sub_694_2_n_111 | (sub_694_2_n_160 & sub_694_2_n_78));
 assign sub_694_2_n_170 = (~sub_694_2_n_5 | (sub_694_2_n_160 & sub_694_2_n_44));
 assign sub_694_2_n_169 = ~(sub_694_2_n_160 & (~sub_694_2_n_121 & ~sub_694_2_n_118));
 assign sub_694_2_n_168 = ~(sub_694_2_n_130 & (sub_694_2_n_159 | sub_694_2_n_121));
 assign n_2294 = ~((sub_694_2_n_159 & ~sub_694_2_n_96) | (sub_694_2_n_160 & sub_694_2_n_96));
 assign sub_694_2_n_166 = ~(sub_694_2_n_112 | (sub_694_2_n_157 & sub_694_2_n_79));
 assign sub_694_2_n_165 = (~sub_694_2_n_14 | (sub_694_2_n_157 & sub_694_2_n_6));
 assign sub_694_2_n_164 = ~(sub_694_2_n_47 & (sub_694_2_n_156 | sub_694_2_n_52));
 assign n_2298 = ~(sub_694_2_n_94 ^ sub_694_2_n_157);
 assign n_2300 = ~(sub_694_2_n_93 ^ sub_694_2_n_156);
 assign n_2301 = ~(sub_694_2_n_91 ^ sub_694_2_n_155);
 assign sub_694_2_n_159 = ~sub_694_2_n_160;
 assign sub_694_2_n_160 = ~(~sub_694_2_n_135 & sub_694_2_n_158);
 assign sub_694_2_n_158 = ~(sub_694_2_n_152 & (~sub_694_2_n_117 & ~sub_694_2_n_120));
 assign sub_694_2_n_157 = ~(sub_694_2_n_128 & (sub_694_2_n_151 | sub_694_2_n_117));
 assign sub_694_2_n_156 = ~(sub_694_2_n_109 | (sub_694_2_n_152 & sub_694_2_n_104));
 assign sub_694_2_n_155 = ~(sub_694_2_n_50 & (sub_694_2_n_151 | sub_694_2_n_17));
 assign n_2302 = ~((sub_694_2_n_151 & ~sub_694_2_n_66) | (sub_694_2_n_152 & sub_694_2_n_66));
 assign n_2303 = ~(sub_694_2_n_76 ^ sub_694_2_n_150);
 assign sub_694_2_n_151 = ~sub_694_2_n_152;
 assign sub_694_2_n_152 = ~(sub_694_2_n_145 & (~sub_694_2_n_36 & ~n_3688));
 assign sub_694_2_n_150 = ~(sub_694_2_n_51 & (sub_694_2_n_147 | sub_694_2_n_22));
 assign n_2304 = (sub_694_2_n_73 ^ sub_694_2_n_147);
 assign n_2305 = (sub_694_2_n_69 ^ sub_694_2_n_146);
 assign sub_694_2_n_147 = ~(sub_694_2_n_115 | (sub_694_2_n_142 & sub_694_2_n_83));
 assign sub_694_2_n_146 = (~sub_694_2_n_3 | (sub_694_2_n_142 & sub_694_2_n_0));
 assign sub_694_2_n_145 = ~(sub_694_2_n_142 & (~sub_694_2_n_106 & ~sub_694_2_n_82));
 assign n_2306 = ~(sub_694_2_n_90 ^ sub_694_2_n_142);
 assign sub_694_2_n_143 = ~(n_3687 & (sub_694_2_n_100 | n_587));
 assign sub_694_2_n_142 = ~(~sub_694_2_n_33 & sub_694_2_n_138);
 assign n_2307 = (sub_694_2_n_88 ^ sub_694_2_n_137);
 assign sub_694_2_n_138 = ~(sub_694_2_n_55 & (sub_694_2_n_19 | (sub_694_2_n_132 & sub_694_2_n_29)));
 assign sub_694_2_n_137 = (sub_694_2_n_19 | (sub_694_2_n_132 & sub_694_2_n_29));
 assign sub_694_2_n_136 = ~(sub_694_2_n_133 | sub_694_2_n_127);
 assign sub_694_2_n_135 = ~(sub_694_2_n_35 & (sub_694_2_n_126 & (sub_694_2_n_128 | sub_694_2_n_120)));
 assign n_2308 = ~(sub_694_2_n_132 ^ sub_694_2_n_74);
 assign sub_694_2_n_133 = ~(sub_694_2_n_61 & (sub_694_2_n_130 | sub_694_2_n_118));
 assign sub_694_2_n_132 = ((sub_694_2_n_13 & n_516) | (n_3517 & (sub_694_2_n_13 ^ n_516)));
 assign n_2309 = (n_3517 ^ (sub_694_2_n_13 ^ n_516));
 assign sub_694_2_n_130 = ~(sub_694_2_n_108 | (sub_694_2_n_111 & sub_694_2_n_80));
 assign sub_694_2_n_129 = ~(sub_694_2_n_107 | (sub_694_2_n_110 & sub_694_2_n_81));
 assign sub_694_2_n_128 = ~(sub_694_2_n_116 | (sub_694_2_n_109 & sub_694_2_n_105));
 assign sub_694_2_n_127 = ~(sub_694_2_n_123 & (sub_694_2_n_53 | sub_694_2_n_31));
 assign sub_694_2_n_126 = ~((~sub_694_2_n_15 & ~sub_694_2_n_27) | (sub_694_2_n_112 & sub_694_2_n_84));
 assign sub_694_2_n_124 = (sub_694_2_n_122 | sub_694_2_n_119);
 assign sub_694_2_n_123 = ~(sub_694_2_n_113 & sub_694_2_n_85);
 assign sub_694_2_n_116 = ~(sub_694_2_n_63 & (sub_694_2_n_47 | sub_694_2_n_46));
 assign sub_694_2_n_122 = ~(sub_694_2_n_102 & sub_694_2_n_81);
 assign sub_694_2_n_121 = ~(sub_694_2_n_78 & sub_694_2_n_80);
 assign sub_694_2_n_120 = ~(sub_694_2_n_79 & sub_694_2_n_84);
 assign sub_694_2_n_119 = ~(~n_587 & (sub_694_2_n_60 & sub_694_2_n_56));
 assign sub_694_2_n_118 = ~(sub_694_2_n_103 & sub_694_2_n_85);
 assign sub_694_2_n_117 = ~(sub_694_2_n_104 & sub_694_2_n_105);
 assign sub_694_2_n_115 = ~sub_694_2_n_114;
 assign sub_694_2_n_108 = ~(sub_694_2_n_58 & (sub_694_2_n_1 | sub_694_2_n_41));
 assign sub_694_2_n_107 = ~(sub_694_2_n_37 & (sub_694_2_n_28 | sub_694_2_n_16));
 assign sub_694_2_n_114 = (~sub_694_2_n_2 & (sub_694_2_n_3 | sub_694_2_n_42));
 assign sub_694_2_n_113 = ~(sub_694_2_n_38 & (sub_694_2_n_24 | sub_694_2_n_32));
 assign sub_694_2_n_112 = ~(sub_694_2_n_54 & (sub_694_2_n_14 | sub_694_2_n_25));
 assign sub_694_2_n_111 = ~(sub_694_2_n_62 & (sub_694_2_n_5 | sub_694_2_n_45));
 assign sub_694_2_n_110 = ~(sub_694_2_n_57 & (sub_694_2_n_43 | sub_694_2_n_20));
 assign sub_694_2_n_109 = ~(sub_694_2_n_59 & (sub_694_2_n_50 | sub_694_2_n_18));
 assign sub_694_2_n_100 = ~(sub_694_2_n_60 & sub_694_2_n_34);
 assign sub_694_2_n_99 = ~(~sub_694_2_n_25 & sub_694_2_n_54);
 assign sub_694_2_n_106 = ~(sub_694_2_n_49 & ~sub_694_2_n_22);
 assign sub_694_2_n_98 = ~(sub_694_2_n_28 & ~sub_694_2_n_26);
 assign sub_694_2_n_97 = ~(~sub_694_2_n_45 & sub_694_2_n_62);
 assign sub_694_2_n_105 = ~(sub_694_2_n_52 | sub_694_2_n_46);
 assign sub_694_2_n_96 = (sub_694_2_n_5 & sub_694_2_n_44);
 assign sub_694_2_n_95 = ~(~sub_694_2_n_15 | sub_694_2_n_23);
 assign sub_694_2_n_94 = ~(sub_694_2_n_14 & sub_694_2_n_6);
 assign sub_694_2_n_104 = ~(sub_694_2_n_17 | sub_694_2_n_18);
 assign sub_694_2_n_93 = ~(~sub_694_2_n_47 | sub_694_2_n_52);
 assign sub_694_2_n_92 = ~(~sub_694_2_n_27 & sub_694_2_n_35);
 assign sub_694_2_n_91 = ~(~sub_694_2_n_18 & sub_694_2_n_59);
 assign sub_694_2_n_103 = ~(~sub_694_2_n_4 | sub_694_2_n_32);
 assign sub_694_2_n_102 = ~(sub_694_2_n_21 | sub_694_2_n_20);
 assign sub_694_2_n_90 = ~(sub_694_2_n_3 & sub_694_2_n_0);
 assign sub_694_2_n_89 = ~(~sub_694_2_n_46 & sub_694_2_n_63);
 assign sub_694_2_n_88 = ~(sub_694_2_n_33 | ~sub_694_2_n_55);
 assign sub_694_2_n_87 = ~(sub_694_2_n_20 | ~sub_694_2_n_57);
 assign sub_694_2_n_86 = ~(~sub_694_2_n_41 & sub_694_2_n_58);
 assign sub_694_2_n_83 = ~sub_694_2_n_82;
 assign n_2310 = ~(sub_694_2_n_39 & (~{in2[3]} | {in1[0]}));
 assign sub_694_2_n_76 = ~(~sub_694_2_n_36 & sub_694_2_n_49);
 assign sub_694_2_n_75 = ~(sub_694_2_n_16 | ~sub_694_2_n_37);
 assign sub_694_2_n_74 = ~(sub_694_2_n_29 & ~sub_694_2_n_19);
 assign sub_694_2_n_85 = ~(sub_694_2_n_30 | sub_694_2_n_31);
 assign sub_694_2_n_73 = ~(sub_694_2_n_51 & ~sub_694_2_n_22);
 assign sub_694_2_n_84 = ~(sub_694_2_n_23 | sub_694_2_n_27);
 assign sub_694_2_n_82 = ~(~sub_694_2_n_42 & sub_694_2_n_0);
 assign sub_694_2_n_72 = ~(~sub_694_2_n_1 | sub_694_2_n_40);
 assign sub_694_2_n_81 = ~(sub_694_2_n_26 | sub_694_2_n_16);
 assign sub_694_2_n_80 = ~(sub_694_2_n_40 | sub_694_2_n_41);
 assign sub_694_2_n_71 = ~(sub_694_2_n_43 & ~sub_694_2_n_21);
 assign sub_694_2_n_70 = ~(sub_694_2_n_31 | ~sub_694_2_n_61);
 assign sub_694_2_n_69 = ~(sub_694_2_n_2 | sub_694_2_n_42);
 assign sub_694_2_n_68 = ~(sub_694_2_n_30 | ~sub_694_2_n_53);
 assign sub_694_2_n_79 = ~(sub_694_2_n_25 | ~sub_694_2_n_6);
 assign sub_694_2_n_67 = ~(sub_694_2_n_38 & ~sub_694_2_n_32);
 assign sub_694_2_n_66 = ~(~sub_694_2_n_50 | sub_694_2_n_17);
 assign sub_694_2_n_65 = ~(sub_694_2_n_24 & sub_694_2_n_4);
 assign sub_694_2_n_78 = ~(sub_694_2_n_45 | ~sub_694_2_n_44);
 assign sub_694_2_n_64 = ~(sub_694_2_n_34 | ~sub_694_2_n_56);
 assign sub_694_2_n_49 = ~sub_694_2_n_48;
 assign sub_694_2_n_63 = ~(~n_428 & n_3523);
 assign sub_694_2_n_62 = ~(~n_561 & n_3530);
 assign sub_694_2_n_61 = ~(~n_459 & n_2258);
 assign sub_694_2_n_60 = ~(n_408 | n_500);
 assign sub_694_2_n_59 = ~(~n_394 & n_3526);
 assign sub_694_2_n_58 = ~(~n_449 & n_3515);
 assign sub_694_2_n_57 = ~(~n_541 & n_2256);
 assign sub_694_2_n_56 = ~(~n_3524 & n_621);
 assign sub_694_2_n_55 = ~(sub_694_2_n_10 & n_531);
 assign sub_694_2_n_54 = ~(~n_348 & n_3519);
 assign sub_694_2_n_53 = ~(~n_337 & n_2259);
 assign sub_694_2_n_52 = ~(~n_358 | n_3535);
 assign sub_694_2_n_51 = ~(~n_653 & n_3531);
 assign sub_694_2_n_50 = ~(sub_694_2_n_12 & n_3527);
 assign sub_694_2_n_48 = ~(~n_676 | n_3529);
 assign sub_694_2_n_47 = ~(~n_358 & n_3535);
 assign sub_694_2_n_46 = ~(~n_428 | n_3523);
 assign sub_694_2_n_45 = ~(~n_561 | n_3530);
 assign sub_694_2_n_44 = ~(~n_3533 & n_469);
 assign sub_694_2_n_43 = ~(sub_694_2_n_9 & n_3520);
 assign sub_694_2_n_42 = ~(~n_635 | n_3532);
 assign sub_694_2_n_41 = ~(~n_449 | n_3515);
 assign sub_694_2_n_40 = ~(~n_607 | n_3528);
 assign sub_694_2_n_39 = ~({in1[0]} & ~{in2[3]});
 assign sub_694_2_n_38 = ~(~n_597 & n_2260);
 assign sub_694_2_n_37 = ~(~n_551 & n_2254);
 assign sub_694_2_n_36 = ~(~n_3529 | n_676);
 assign sub_694_2_n_35 = ~(~n_520 & n_3516);
 assign sub_694_2_n_34 = ~(~n_3524 | n_621);
 assign sub_694_2_n_33 = ~(n_531 | sub_694_2_n_10);
 assign sub_694_2_n_32 = ~(~n_597 | n_2260);
 assign sub_694_2_n_31 = ~(~n_459 | n_2258);
 assign sub_694_2_n_30 = ~(~n_337 | n_2259);
 assign sub_694_2_n_29 = ~(sub_694_2_n_11 & n_418);
 assign sub_694_2_n_28 = ~(~n_663 & n_2255);
 assign sub_694_2_n_27 = ~(~n_520 | n_3516);
 assign sub_694_2_n_26 = ~(~n_663 | n_2255);
 assign sub_694_2_n_25 = ~(~n_348 | n_3519);
 assign sub_694_2_n_24 = ~(~n_479 & n_3521);
 assign sub_694_2_n_23 = ~(~n_369 | n_3518);
 assign sub_694_2_n_22 = ~(~n_653 | n_3531);
 assign sub_694_2_n_21 = ~(n_3520 | sub_694_2_n_9);
 assign sub_694_2_n_20 = ~(~n_541 | n_2256);
 assign sub_694_2_n_19 = ~(n_418 | sub_694_2_n_11);
 assign sub_694_2_n_18 = ~(~n_394 | n_3526);
 assign sub_694_2_n_17 = ~(n_3527 | sub_694_2_n_12);
 assign sub_694_2_n_16 = ~(~n_551 | n_2254);
 assign sub_694_2_n_15 = ~(~n_369 & n_3518);
 assign sub_694_2_n_14 = ~(~n_686 & n_3522);
 assign sub_694_2_n_13 = ~n_384;
 assign sub_694_2_n_12 = ~n_438;
 assign sub_694_2_n_11 = ~n_3068;
 assign sub_694_2_n_10 = ~n_3525;
 assign sub_694_2_n_9 = ~n_1108;
 assign sub_694_2_n_6 = ~(~n_3522 & n_686);
 assign sub_694_2_n_5 = ~(~n_469 & n_3533);
 assign sub_694_2_n_4 = ~(~n_3521 & n_479);
 assign sub_694_2_n_3 = ~(~n_698 & n_3534);
 assign sub_694_2_n_2 = ~(n_635 | ~n_3532);
 assign sub_694_2_n_1 = ~(~n_607 & n_3528);
 assign sub_694_2_n_0 = ~(~n_3534 & n_698);
 assign sub_713_2_n_1 = (sub_713_2_n_131 & ~(sub_713_2_n_161 & sub_713_2_n_118));
 assign n_2341 = (sub_713_2_n_76 ^ sub_713_2_n_188);
 assign n_2343 = (sub_713_2_n_72 ^ sub_713_2_n_187);
 assign n_2347 = (sub_713_2_n_66 ^ sub_713_2_n_186);
 assign sub_713_2_n_188 = ~(sub_713_2_n_17 & (sub_713_2_n_1 | sub_713_2_n_49));
 assign sub_713_2_n_187 = ~(sub_713_2_n_14 & (sub_713_2_n_178 | sub_713_2_n_36));
 assign sub_713_2_n_186 = ~(sub_713_2_n_53 & (sub_713_2_n_174 | sub_713_2_n_12));
 assign n_2349 = (sub_713_2_n_92 ^ sub_713_2_n_176);
 assign n_2351 = ~(sub_713_2_n_98 ^ sub_713_2_n_175);
 assign n_2342 = (sub_713_2_n_74 ^ sub_713_2_n_1);
 assign n_2344 = (sub_713_2_n_70 ^ sub_713_2_n_178);
 assign n_2345 = (sub_713_2_n_69 ^ sub_713_2_n_169);
 assign n_2348 = (sub_713_2_n_99 ^ sub_713_2_n_174);
 assign n_2355 = ~(sub_713_2_n_89 ^ sub_713_2_n_167);
 assign n_2340 = (sub_713_2_n_121 & (sub_713_2_n_168 & (sub_713_2_n_131 | sub_713_2_n_115)));
 assign sub_713_2_n_176 = ~(sub_713_2_n_45 & (sub_713_2_n_160 | sub_713_2_n_40));
 assign sub_713_2_n_175 = ~(sub_713_2_n_10 & (sub_713_2_n_163 | sub_713_2_n_15));
 assign sub_713_2_n_178 = ~(sub_713_2_n_114 | (sub_713_2_n_161 & sub_713_2_n_82));
 assign n_2352 = ~(sub_713_2_n_95 ^ sub_713_2_n_163);
 assign n_2350 = ~(sub_713_2_n_101 ^ sub_713_2_n_160);
 assign n_2346 = (sub_713_2_n_67 ^ sub_713_2_n_161);
 assign n_2353 = ~(sub_713_2_n_94 ^ sub_713_2_n_162);
 assign sub_713_2_n_169 = (~sub_713_2_n_6 | (sub_713_2_n_161 & sub_713_2_n_21));
 assign sub_713_2_n_174 = (~sub_713_2_n_109 & (sub_713_2_n_160 | sub_713_2_n_106));
 assign sub_713_2_n_168 = ~(sub_713_2_n_125 & (sub_713_2_n_136 | (sub_713_2_n_152 & sub_713_2_n_123)));
 assign sub_713_2_n_167 = ~(sub_713_2_n_16 & (sub_713_2_n_158 | sub_713_2_n_19));
 assign n_2356 = ~(sub_713_2_n_91 ^ sub_713_2_n_158);
 assign n_2357 = ~(sub_713_2_n_88 ^ sub_713_2_n_157);
 assign n_2359 = ~(sub_713_2_n_65 ^ sub_713_2_n_156);
 assign sub_713_2_n_163 = ~(sub_713_2_n_111 | (sub_713_2_n_152 & sub_713_2_n_83));
 assign sub_713_2_n_162 = (~sub_713_2_n_5 | (sub_713_2_n_152 & sub_713_2_n_39));
 assign sub_713_2_n_161 = (sub_713_2_n_136 | (sub_713_2_n_152 & sub_713_2_n_123));
 assign sub_713_2_n_160 = ~(sub_713_2_n_132 | (sub_713_2_n_152 & sub_713_2_n_117));
 assign n_2354 = ~(sub_713_2_n_93 ^ sub_713_2_n_152);
 assign sub_713_2_n_158 = ~(sub_713_2_n_110 | (sub_713_2_n_151 & sub_713_2_n_104));
 assign sub_713_2_n_157 = (~sub_713_2_n_8 | (sub_713_2_n_151 & sub_713_2_n_50));
 assign sub_713_2_n_156 = ~(sub_713_2_n_41 & (sub_713_2_n_150 | sub_713_2_n_48));
 assign n_2358 = ~(sub_713_2_n_90 ^ sub_713_2_n_151);
 assign n_2360 = ~(sub_713_2_n_96 ^ sub_713_2_n_150);
 assign n_2361 = ~(sub_713_2_n_100 ^ sub_713_2_n_149);
 assign sub_713_2_n_152 = ~(sub_713_2_n_135 & (sub_713_2_n_146 | (sub_713_2_n_119 | sub_713_2_n_116)));
 assign sub_713_2_n_151 = ~(sub_713_2_n_133 & (sub_713_2_n_146 | sub_713_2_n_119));
 assign sub_713_2_n_150 = (~sub_713_2_n_113 & (sub_713_2_n_146 | sub_713_2_n_86));
 assign sub_713_2_n_149 = ~(sub_713_2_n_38 & (sub_713_2_n_146 | sub_713_2_n_54));
 assign n_2362 = ~(sub_713_2_n_68 ^ sub_713_2_n_146);
 assign n_2363 = ~(sub_713_2_n_0 ^ sub_713_2_n_145);
 assign sub_713_2_n_146 = ~(sub_713_2_n_140 | (sub_713_2_n_27 | sub_713_2_n_128));
 assign sub_713_2_n_145 = ~(sub_713_2_n_43 | (sub_713_2_n_142 & sub_713_2_n_47));
 assign n_2364 = (sub_713_2_n_71 ^ sub_713_2_n_142);
 assign n_2365 = (sub_713_2_n_64 ^ sub_713_2_n_141);
 assign sub_713_2_n_142 = ~(sub_713_2_n_112 & (sub_713_2_n_138 | sub_713_2_n_80));
 assign sub_713_2_n_141 = ~(sub_713_2_n_20 & (sub_713_2_n_138 | sub_713_2_n_7));
 assign sub_713_2_n_140 = ~(sub_713_2_n_138 | (sub_713_2_n_80 | sub_713_2_n_105));
 assign n_2366 = (sub_713_2_n_75 ^ sub_713_2_n_138);
 assign sub_713_2_n_138 = ~(sub_713_2_n_63 | (sub_713_2_n_2 & sub_713_2_n_55));
 assign n_2367 = (sub_713_2_n_97 ^ sub_713_2_n_2);
 assign sub_713_2_n_136 = (sub_713_2_n_57 | (sub_713_2_n_130 | (sub_713_2_n_132 & sub_713_2_n_120)));
 assign sub_713_2_n_135 = (sub_713_2_n_31 & (sub_713_2_n_129 & (sub_713_2_n_133 | sub_713_2_n_116)));
 assign n_2368 = (sub_713_2_n_127 ^ sub_713_2_n_87);
 assign sub_713_2_n_133 = ~(sub_713_2_n_103 | (sub_713_2_n_62 | (sub_713_2_n_113 & sub_713_2_n_107)));
 assign sub_713_2_n_132 = ~(sub_713_2_n_26 & (sub_713_2_n_124 & (sub_713_2_n_10 | sub_713_2_n_42)));
 assign sub_713_2_n_131 = ~(sub_713_2_n_77 | (sub_713_2_n_29 | (sub_713_2_n_114 & sub_713_2_n_81)));
 assign sub_713_2_n_130 = ~(sub_713_2_n_122 & (sub_713_2_n_53 | sub_713_2_n_18));
 assign sub_713_2_n_129 = ~((~sub_713_2_n_16 & ~sub_713_2_n_44) | (sub_713_2_n_110 & sub_713_2_n_85));
 assign sub_713_2_n_128 = ~(sub_713_2_n_102 & (sub_713_2_n_112 | sub_713_2_n_105));
 assign sub_713_2_n_127 = ~(sub_713_2_n_25 | (n_509 & sub_713_2_n_33));
 assign n_2369 = (n_509 ^ sub_713_2_n_73);
 assign sub_713_2_n_125 = ~(sub_713_2_n_115 | ~sub_713_2_n_118);
 assign sub_713_2_n_124 = ~(sub_713_2_n_111 & sub_713_2_n_108);
 assign sub_713_2_n_123 = (sub_713_2_n_117 & sub_713_2_n_120);
 assign sub_713_2_n_122 = ~(sub_713_2_n_109 & sub_713_2_n_84);
 assign sub_713_2_n_121 = ~(sub_713_2_n_60 & (sub_713_2_n_78 | sub_713_2_n_61));
 assign sub_713_2_n_120 = ~(~sub_713_2_n_84 | sub_713_2_n_106);
 assign sub_713_2_n_119 = ~(~sub_713_2_n_86 & sub_713_2_n_107);
 assign sub_713_2_n_118 = (sub_713_2_n_82 & sub_713_2_n_81);
 assign sub_713_2_n_117 = (sub_713_2_n_83 & sub_713_2_n_108);
 assign sub_713_2_n_116 = ~(sub_713_2_n_104 & sub_713_2_n_85);
 assign sub_713_2_n_115 = ~(~sub_713_2_n_49 & (sub_713_2_n_22 & sub_713_2_n_60));
 assign sub_713_2_n_114 = ~(sub_713_2_n_59 & (sub_713_2_n_6 | sub_713_2_n_46));
 assign sub_713_2_n_113 = ~(sub_713_2_n_56 & (sub_713_2_n_38 | sub_713_2_n_52));
 assign sub_713_2_n_112 = (~sub_713_2_n_58 & (sub_713_2_n_20 | sub_713_2_n_11));
 assign sub_713_2_n_111 = ~(sub_713_2_n_28 & (sub_713_2_n_5 | sub_713_2_n_13));
 assign sub_713_2_n_110 = ~(sub_713_2_n_32 & (sub_713_2_n_8 | sub_713_2_n_9));
 assign sub_713_2_n_109 = ~(sub_713_2_n_30 & (sub_713_2_n_45 | sub_713_2_n_35));
 assign sub_713_2_n_103 = ~(sub_713_2_n_41 | sub_713_2_n_37);
 assign sub_713_2_n_102 = ~(sub_713_2_n_43 & sub_713_2_n_51);
 assign sub_713_2_n_101 = ~(~sub_713_2_n_45 | sub_713_2_n_40);
 assign sub_713_2_n_108 = ~(sub_713_2_n_15 | sub_713_2_n_42);
 assign sub_713_2_n_100 = ~(~sub_713_2_n_52 & sub_713_2_n_56);
 assign sub_713_2_n_99 = ~(sub_713_2_n_53 & ~sub_713_2_n_12);
 assign sub_713_2_n_98 = ~(sub_713_2_n_26 & ~sub_713_2_n_42);
 assign sub_713_2_n_97 = ~(sub_713_2_n_63 | ~sub_713_2_n_55);
 assign sub_713_2_n_96 = ~(~sub_713_2_n_41 | sub_713_2_n_48);
 assign sub_713_2_n_95 = ~(~sub_713_2_n_10 | sub_713_2_n_15);
 assign sub_713_2_n_94 = ~(~sub_713_2_n_13 & sub_713_2_n_28);
 assign sub_713_2_n_107 = ~(sub_713_2_n_48 | sub_713_2_n_37);
 assign sub_713_2_n_93 = ~(sub_713_2_n_5 & sub_713_2_n_39);
 assign sub_713_2_n_106 = (sub_713_2_n_40 | sub_713_2_n_35);
 assign sub_713_2_n_92 = ~(sub_713_2_n_35 | ~sub_713_2_n_30);
 assign sub_713_2_n_91 = ~(~sub_713_2_n_16 | sub_713_2_n_19);
 assign sub_713_2_n_90 = ~(sub_713_2_n_8 & sub_713_2_n_50);
 assign sub_713_2_n_89 = ~(sub_713_2_n_31 & ~sub_713_2_n_44);
 assign sub_713_2_n_88 = ~(~sub_713_2_n_9 & sub_713_2_n_32);
 assign sub_713_2_n_105 = ~(sub_713_2_n_47 & sub_713_2_n_51);
 assign sub_713_2_n_87 = ~(sub_713_2_n_34 & ~sub_713_2_n_23);
 assign sub_713_2_n_104 = ~(~sub_713_2_n_50 | sub_713_2_n_9);
 assign n_2370 = ~(sub_713_2_n_4 & (~{in2[2]} | {in1[0]}));
 assign sub_713_2_n_78 = ~(~sub_713_2_n_22 | sub_713_2_n_17);
 assign sub_713_2_n_77 = ~(sub_713_2_n_14 | sub_713_2_n_24);
 assign sub_713_2_n_86 = (sub_713_2_n_54 | sub_713_2_n_52);
 assign sub_713_2_n_76 = ~(sub_713_2_n_61 | ~sub_713_2_n_22);
 assign sub_713_2_n_75 = ~(~sub_713_2_n_7 & sub_713_2_n_20);
 assign sub_713_2_n_74 = ~(sub_713_2_n_17 & ~sub_713_2_n_49);
 assign sub_713_2_n_73 = ~(sub_713_2_n_25 | ~sub_713_2_n_33);
 assign sub_713_2_n_72 = ~(sub_713_2_n_29 | sub_713_2_n_24);
 assign sub_713_2_n_85 = ~(sub_713_2_n_19 | sub_713_2_n_44);
 assign sub_713_2_n_71 = ~(sub_713_2_n_43 | ~sub_713_2_n_47);
 assign sub_713_2_n_70 = ~(sub_713_2_n_14 & ~sub_713_2_n_36);
 assign sub_713_2_n_84 = ~(sub_713_2_n_12 | sub_713_2_n_18);
 assign sub_713_2_n_69 = ~(sub_713_2_n_46 | ~sub_713_2_n_59);
 assign sub_713_2_n_83 = ~(sub_713_2_n_13 | ~sub_713_2_n_39);
 assign sub_713_2_n_68 = ~(~sub_713_2_n_38 | sub_713_2_n_54);
 assign sub_713_2_n_67 = (sub_713_2_n_6 & sub_713_2_n_21);
 assign sub_713_2_n_82 = ~(sub_713_2_n_46 | ~sub_713_2_n_21);
 assign sub_713_2_n_66 = ~(sub_713_2_n_57 | sub_713_2_n_18);
 assign sub_713_2_n_81 = ~(sub_713_2_n_36 | sub_713_2_n_24);
 assign sub_713_2_n_65 = (sub_713_2_n_62 | sub_713_2_n_37);
 assign sub_713_2_n_64 = ~(sub_713_2_n_58 | sub_713_2_n_11);
 assign sub_713_2_n_80 = (sub_713_2_n_7 | sub_713_2_n_11);
 assign sub_713_2_n_63 = ~(~n_1021 | n_530);
 assign sub_713_2_n_62 = ~(~n_1036 | n_427);
 assign sub_713_2_n_61 = ~(~n_1032 | n_586);
 assign sub_713_2_n_60 = ~(n_407 | n_499);
 assign sub_713_2_n_59 = ~(~n_540 & n_1030);
 assign sub_713_2_n_58 = ~(~n_1042 | n_634);
 assign sub_713_2_n_57 = ~(~n_1020 | n_458);
 assign sub_713_2_n_56 = ~(~n_393 & n_1033);
 assign sub_713_2_n_55 = ~(~n_1021 & n_530);
 assign sub_713_2_n_54 = ~(~n_437 | n_1040);
 assign sub_713_2_n_53 = ~(~n_336 & n_1019);
 assign sub_713_2_n_52 = ~(~n_393 | n_1033);
 assign sub_713_2_n_51 = ~(~n_1039 & n_675);
 assign sub_713_2_n_50 = ~(~n_1023 & n_685);
 assign sub_713_2_n_49 = ~(~n_620 | n_2312);
 assign sub_713_2_n_48 = ~(~n_357 | n_1034);
 assign sub_713_2_n_47 = ~(~n_1041 & n_652);
 assign sub_713_2_n_46 = ~(~n_540 | n_1030);
 assign sub_713_2_n_45 = ~(~n_478 & n_1037);
 assign sub_713_2_n_44 = ~(~n_519 | n_1028);
 assign sub_713_2_n_43 = ~(~n_1041 | n_652);
 assign sub_713_2_n_42 = ~(~n_448 | n_1027);
 assign sub_713_2_n_41 = ~(~n_357 & n_1034);
 assign sub_713_2_n_40 = ~(~n_478 | n_1037);
 assign sub_713_2_n_39 = ~(n_468 & ~n_1017);
 assign sub_713_2_n_38 = ~(~n_437 & n_1040);
 assign sub_713_2_n_37 = ~(~n_427 | n_1036);
 assign sub_713_2_n_36 = ~(~n_662 | n_1022);
 assign sub_713_2_n_35 = ~(~n_596 | n_1035);
 assign sub_713_2_n_34 = ~(~n_417 & n_1025);
 assign sub_713_2_n_33 = ~(~n_1026 & n_383);
 assign sub_713_2_n_32 = ~(~n_347 & n_1031);
 assign sub_713_2_n_31 = ~(~n_519 & n_1028);
 assign sub_713_2_n_30 = ~(~n_596 & n_1035);
 assign sub_713_2_n_29 = ~(~n_1018 | n_550);
 assign sub_713_2_n_28 = ~(~n_560 & n_1043);
 assign sub_713_2_n_27 = ~(~n_1039 | n_675);
 assign sub_713_2_n_26 = ~(~n_448 & n_1027);
 assign sub_713_2_n_25 = ~(~n_1026 | n_383);
 assign sub_713_2_n_24 = ~(~n_550 | n_1018);
 assign sub_713_2_n_23 = ~(~n_417 | n_1025);
 assign sub_713_2_n_22 = ~(n_586 & ~n_1032);
 assign sub_713_2_n_21 = ~(n_1107 & ~n_1016);
 assign sub_713_2_n_20 = ~(~n_697 & n_1044);
 assign sub_713_2_n_19 = ~(~n_368 | n_1029);
 assign sub_713_2_n_18 = ~(~n_458 | n_1020);
 assign sub_713_2_n_17 = ~(~n_620 & n_2312);
 assign sub_713_2_n_16 = ~(~n_368 & n_1029);
 assign sub_713_2_n_15 = ~(~n_606 | n_1038);
 assign sub_713_2_n_14 = ~(~n_662 & n_1022);
 assign sub_713_2_n_13 = ~(~n_560 | n_1043);
 assign sub_713_2_n_12 = ~(~n_336 | n_1019);
 assign sub_713_2_n_11 = ~(~n_634 | n_1042);
 assign sub_713_2_n_10 = ~(~n_606 & n_1038);
 assign sub_713_2_n_9 = ~(~n_347 | n_1031);
 assign sub_713_2_n_8 = ~(~n_685 & n_1023);
 assign sub_713_2_n_7 = ~(~n_697 | n_1044);
 assign sub_713_2_n_6 = ~(~n_1107 & n_1016);
 assign sub_713_2_n_5 = ~(~n_468 & n_1017);
 assign sub_713_2_n_4 = ~({in1[0]} & ~{in2[2]});
 assign sub_713_2_n_2 = ~(sub_713_2_n_34 & (sub_713_2_n_127 | sub_713_2_n_23));
 assign sub_713_2_n_0 = ~(sub_713_2_n_27 | ~sub_713_2_n_51);
 assign sub_732_2_n_1 = (sub_732_2_n_133 & ~(sub_732_2_n_164 & sub_732_2_n_118));
 assign n_2402 = ~(sub_732_2_n_75 ^ sub_732_2_n_193);
 assign n_2403 = ~(sub_732_2_n_74 ^ sub_732_2_n_192);
 assign n_2405 = ~(sub_732_2_n_69 ^ sub_732_2_n_191);
 assign n_2409 = ~(sub_732_2_n_64 ^ sub_732_2_n_194);
 assign sub_732_2_n_194 = ~(sub_732_2_n_5 & (sub_732_2_n_183 | n_1065));
 assign sub_732_2_n_193 = ~(sub_732_2_n_110 & (sub_732_2_n_1 | sub_732_2_n_83));
 assign sub_732_2_n_192 = ~(sub_732_2_n_42 & (sub_732_2_n_1 | sub_732_2_n_50));
 assign sub_732_2_n_191 = ~(sub_732_2_n_38 & (sub_732_2_n_179 | sub_732_2_n_48));
 assign n_2410 = (sub_732_2_n_101 ^ sub_732_2_n_183);
 assign n_2411 = ~(sub_732_2_n_100 ^ sub_732_2_n_180);
 assign n_2413 = (sub_732_2_n_97 ^ sub_732_2_n_181);
 assign n_2404 = ~(sub_732_2_n_73 ^ sub_732_2_n_1);
 assign n_2406 = ~(sub_732_2_n_68 ^ sub_732_2_n_179);
 assign n_2407 = ~(sub_732_2_n_66 ^ sub_732_2_n_174);
 assign n_2417 = (n_1055 ^ n_1091);
 assign n_2401 = (sub_732_2_n_132 & (sub_732_2_n_173 & (sub_732_2_n_133 | sub_732_2_n_121)));
 assign sub_732_2_n_181 = ~(sub_732_2_n_41 & (sub_732_2_n_166 | n_1101));
 assign sub_732_2_n_180 = ~(n_1056 & (sub_732_2_n_168 | n_1057));
 assign sub_732_2_n_183 = ~(sub_732_2_n_109 | (sub_732_2_n_167 & sub_732_2_n_105));
 assign n_2414 = (sub_732_2_n_93 ^ sub_732_2_n_166);
 assign n_2412 = ~((sub_732_2_n_168 & ~sub_732_2_n_67) | (sub_732_2_n_167 & sub_732_2_n_67));
 assign n_2408 = ~(sub_732_2_n_76 ^ sub_732_2_n_164);
 assign n_2415 = (sub_732_2_n_92 ^ sub_732_2_n_165);
 assign sub_732_2_n_174 = (~sub_732_2_n_46 | (sub_732_2_n_164 & sub_732_2_n_17));
 assign sub_732_2_n_179 = ~(sub_732_2_n_114 | (sub_732_2_n_164 & sub_732_2_n_85));
 assign sub_732_2_n_173 = ~(sub_732_2_n_126 & (sub_732_2_n_139 | (n_1096 & sub_732_2_n_123)));
 assign sub_732_2_n_172 = ~(sub_732_2_n_10 & (sub_732_2_n_162 | sub_732_2_n_7));
 assign n_2418 = ~(sub_732_2_n_95 ^ sub_732_2_n_162);
 assign n_2419 = ~(sub_732_2_n_89 ^ sub_732_2_n_161);
 assign n_2421 = ~(sub_732_2_n_0 ^ sub_732_2_n_160);
 assign sub_732_2_n_167 = ~sub_732_2_n_168;
 assign sub_732_2_n_168 = ~(sub_732_2_n_134 | (n_1096 & sub_732_2_n_117));
 assign sub_732_2_n_166 = ~(sub_732_2_n_111 | (n_1096 & sub_732_2_n_84));
 assign sub_732_2_n_165 = (~n_1061 | (n_1096 & n_1062));
 assign sub_732_2_n_164 = (sub_732_2_n_139 | (n_1096 & sub_732_2_n_123));
 assign n_2416 = (sub_732_2_n_88 ^ n_1096);
 assign sub_732_2_n_162 = ~(sub_732_2_n_115 | (sub_732_2_n_155 & sub_732_2_n_108));
 assign sub_732_2_n_161 = (~sub_732_2_n_19 | (sub_732_2_n_155 & sub_732_2_n_51));
 assign sub_732_2_n_160 = ~(sub_732_2_n_39 & (sub_732_2_n_154 | sub_732_2_n_13));
 assign n_2422 = ~(sub_732_2_n_87 ^ sub_732_2_n_154);
 assign n_2423 = ~(sub_732_2_n_96 ^ sub_732_2_n_153);
 assign n_2420 = ~(sub_732_2_n_65 ^ sub_732_2_n_155);
 assign sub_732_2_n_156 = ~(sub_732_2_n_138 & (sub_732_2_n_150 | (sub_732_2_n_116 | sub_732_2_n_120)));
 assign sub_732_2_n_155 = ~(sub_732_2_n_135 & (sub_732_2_n_150 | sub_732_2_n_116));
 assign sub_732_2_n_154 = (~sub_732_2_n_113 & (sub_732_2_n_150 | sub_732_2_n_104));
 assign sub_732_2_n_153 = ~(sub_732_2_n_44 & (sub_732_2_n_150 | sub_732_2_n_2));
 assign n_2424 = ~(sub_732_2_n_98 ^ sub_732_2_n_150);
 assign n_2425 = ~(sub_732_2_n_71 ^ sub_732_2_n_149);
 assign sub_732_2_n_150 = ~(sub_732_2_n_144 | (sub_732_2_n_23 | sub_732_2_n_131));
 assign sub_732_2_n_149 = ~(sub_732_2_n_4 & (sub_732_2_n_146 | sub_732_2_n_45));
 assign n_2426 = (sub_732_2_n_90 ^ sub_732_2_n_146);
 assign n_2427 = (sub_732_2_n_94 ^ sub_732_2_n_145);
 assign sub_732_2_n_146 = ~(sub_732_2_n_112 | (sub_732_2_n_142 & sub_732_2_n_81));
 assign sub_732_2_n_145 = (~sub_732_2_n_47 | (sub_732_2_n_142 & sub_732_2_n_3));
 assign sub_732_2_n_144 = (sub_732_2_n_142 & (sub_732_2_n_79 & sub_732_2_n_81));
 assign n_2428 = (sub_732_2_n_99 ^ sub_732_2_n_142);
 assign sub_732_2_n_142 = ~(sub_732_2_n_29 & (sub_732_2_n_28 | (sub_732_2_n_136 & sub_732_2_n_20)));
 assign n_2429 = (sub_732_2_n_70 ^ sub_732_2_n_140);
 assign sub_732_2_n_140 = ~(sub_732_2_n_20 & (sub_732_2_n_128 | sub_732_2_n_18));
 assign sub_732_2_n_139 = (sub_732_2_n_27 | (sub_732_2_n_130 | (sub_732_2_n_134 & sub_732_2_n_119)));
 assign sub_732_2_n_138 = (sub_732_2_n_57 & (sub_732_2_n_129 & (sub_732_2_n_135 | sub_732_2_n_120)));
 assign n_2430 = (sub_732_2_n_72 ^ sub_732_2_n_128);
 assign sub_732_2_n_136 = (sub_732_2_n_128 | sub_732_2_n_18);
 assign sub_732_2_n_135 = ~(sub_732_2_n_102 | (sub_732_2_n_62 | (sub_732_2_n_113 & sub_732_2_n_107)));
 assign sub_732_2_n_134 = ~(sub_732_2_n_56 & (sub_732_2_n_124 & (sub_732_2_n_41 | n_1049)));
 assign sub_732_2_n_133 = ~(sub_732_2_n_78 | (sub_732_2_n_24 | (sub_732_2_n_114 & sub_732_2_n_106)));
 assign sub_732_2_n_132 = ((sub_732_2_n_32 | n_498) & (sub_732_2_n_110 | sub_732_2_n_103));
 assign sub_732_2_n_131 = ~(sub_732_2_n_125 & (sub_732_2_n_4 | sub_732_2_n_37));
 assign sub_732_2_n_130 = ~(sub_732_2_n_122 & (sub_732_2_n_5 | n_1054));
 assign sub_732_2_n_129 = ~((~sub_732_2_n_10 & ~sub_732_2_n_53) | (sub_732_2_n_115 & sub_732_2_n_82));
 assign sub_732_2_n_128 = ~(sub_732_2_n_61 | (n_673 & sub_732_2_n_60));
 assign n_2431 = (n_673 ^ sub_732_2_n_63);
 assign sub_732_2_n_126 = ~(sub_732_2_n_121 | ~sub_732_2_n_118);
 assign sub_732_2_n_125 = ~(sub_732_2_n_112 & sub_732_2_n_79);
 assign sub_732_2_n_124 = ~(sub_732_2_n_111 & sub_732_2_n_86);
 assign sub_732_2_n_123 = (sub_732_2_n_117 & sub_732_2_n_119);
 assign sub_732_2_n_122 = ~(sub_732_2_n_109 & sub_732_2_n_80);
 assign sub_732_2_n_121 = (sub_732_2_n_83 | sub_732_2_n_103);
 assign sub_732_2_n_120 = ~(sub_732_2_n_108 & sub_732_2_n_82);
 assign sub_732_2_n_119 = (sub_732_2_n_105 & sub_732_2_n_80);
 assign sub_732_2_n_118 = (sub_732_2_n_85 & sub_732_2_n_106);
 assign sub_732_2_n_117 = (sub_732_2_n_84 & sub_732_2_n_86);
 assign sub_732_2_n_116 = ~(~sub_732_2_n_104 & sub_732_2_n_107);
 assign sub_732_2_n_115 = ~(sub_732_2_n_22 & (sub_732_2_n_19 | sub_732_2_n_12));
 assign sub_732_2_n_114 = ~(sub_732_2_n_58 & (sub_732_2_n_46 | sub_732_2_n_52));
 assign sub_732_2_n_113 = ~(sub_732_2_n_59 & (sub_732_2_n_44 | sub_732_2_n_40));
 assign sub_732_2_n_112 = ~(sub_732_2_n_30 & (sub_732_2_n_47 | sub_732_2_n_9));
 assign sub_732_2_n_111 = ~(n_1051 & (n_1061 | n_1050));
 assign sub_732_2_n_110 = (~sub_732_2_n_26 & (sub_732_2_n_42 | sub_732_2_n_49));
 assign sub_732_2_n_109 = ~(sub_732_2_n_55 & (n_1056 | n_1082));
 assign sub_732_2_n_102 = ~(sub_732_2_n_39 | sub_732_2_n_43);
 assign sub_732_2_n_108 = ~(~sub_732_2_n_51 | sub_732_2_n_12);
 assign sub_732_2_n_101 = ~(sub_732_2_n_5 & ~n_1065);
 assign sub_732_2_n_100 = ~(sub_732_2_n_55 & ~n_1082);
 assign sub_732_2_n_99 = (sub_732_2_n_47 & sub_732_2_n_3);
 assign sub_732_2_n_98 = ~(~sub_732_2_n_44 | sub_732_2_n_2);
 assign sub_732_2_n_97 = ~(n_1049 | ~sub_732_2_n_56);
 assign sub_732_2_n_96 = ~(sub_732_2_n_59 & ~sub_732_2_n_40);
 assign sub_732_2_n_95 = ~(~sub_732_2_n_10 | sub_732_2_n_7);
 assign sub_732_2_n_94 = ~(sub_732_2_n_9 | ~sub_732_2_n_30);
 assign sub_732_2_n_93 = ~(~n_1101 & sub_732_2_n_41);
 assign sub_732_2_n_92 = ~(n_1050 | ~n_1051);
 assign sub_732_2_n_107 = ~(sub_732_2_n_13 | sub_732_2_n_43);
 assign sub_732_2_n_106 = ~(sub_732_2_n_48 | sub_732_2_n_15);
 assign sub_732_2_n_91 = ~(sub_732_2_n_53 | ~sub_732_2_n_57);
 assign sub_732_2_n_90 = ~(~sub_732_2_n_45 & sub_732_2_n_4);
 assign sub_732_2_n_89 = ~(~sub_732_2_n_12 & sub_732_2_n_22);
 assign sub_732_2_n_88 = (n_1061 & n_1062);
 assign sub_732_2_n_105 = ~(n_1057 | n_1082);
 assign sub_732_2_n_104 = (sub_732_2_n_2 | sub_732_2_n_40);
 assign sub_732_2_n_87 = ~(~sub_732_2_n_39 | sub_732_2_n_13);
 assign sub_732_2_n_103 = ~(~n_498 & sub_732_2_n_31);
 assign sub_732_2_n_78 = ~(sub_732_2_n_38 | sub_732_2_n_15);
 assign n_2432 = ~(sub_732_2_n_33 & (~{in2[1]} | {in1[0]}));
 assign sub_732_2_n_76 = ~(sub_732_2_n_46 & sub_732_2_n_17);
 assign sub_732_2_n_86 = ~(n_1101 | n_1049);
 assign sub_732_2_n_85 = ~(sub_732_2_n_52 | ~sub_732_2_n_17);
 assign sub_732_2_n_84 = ~(n_1050 | ~n_1062);
 assign sub_732_2_n_75 = ~(sub_732_2_n_32 & sub_732_2_n_31);
 assign sub_732_2_n_83 = (sub_732_2_n_50 | sub_732_2_n_49);
 assign sub_732_2_n_74 = (sub_732_2_n_26 | sub_732_2_n_49);
 assign sub_732_2_n_73 = ~(~sub_732_2_n_42 | sub_732_2_n_50);
 assign sub_732_2_n_72 = ~(sub_732_2_n_20 & ~sub_732_2_n_18);
 assign sub_732_2_n_71 = (sub_732_2_n_23 | sub_732_2_n_37);
 assign sub_732_2_n_70 = ~(sub_732_2_n_28 | ~sub_732_2_n_29);
 assign sub_732_2_n_69 = (sub_732_2_n_24 | sub_732_2_n_15);
 assign sub_732_2_n_82 = ~(sub_732_2_n_7 | sub_732_2_n_53);
 assign sub_732_2_n_81 = ~(sub_732_2_n_9 | ~sub_732_2_n_3);
 assign sub_732_2_n_68 = ~(~sub_732_2_n_38 | sub_732_2_n_48);
 assign sub_732_2_n_67 = ~(n_1057 | ~n_1056);
 assign sub_732_2_n_66 = ~(~sub_732_2_n_52 & sub_732_2_n_58);
 assign sub_732_2_n_65 = ~(sub_732_2_n_19 & sub_732_2_n_51);
 assign sub_732_2_n_80 = ~(n_1065 | n_1054);
 assign sub_732_2_n_79 = ~(sub_732_2_n_45 | sub_732_2_n_37);
 assign sub_732_2_n_64 = (sub_732_2_n_27 | n_1054);
 assign sub_732_2_n_63 = ~(~sub_732_2_n_60 | sub_732_2_n_61);
 assign sub_732_2_n_62 = ~(~n_2390 | n_427);
 assign sub_732_2_n_61 = ~(n_383 | ~n_2400);
 assign sub_732_2_n_60 = ~(n_383 & ~n_2400);
 assign sub_732_2_n_59 = ~(~n_393 & n_2392);
 assign sub_732_2_n_58 = ~(~n_539 & n_1084);
 assign sub_732_2_n_57 = ~(~n_519 & n_2386);
 assign sub_732_2_n_56 = ~(~n_447 & n_1052);
 assign sub_732_2_n_55 = ~(~n_595 & n_1085);
 assign sub_732_2_n_54 = ~(~n_596 | n_2380);
 assign sub_732_2_n_53 = ~(~n_519 | n_2386);
 assign sub_732_2_n_52 = ~(~n_539 | n_1084);
 assign sub_732_2_n_51 = ~(~n_2389 & n_685);
 assign sub_732_2_n_50 = ~(~n_619 | n_1081);
 assign sub_732_2_n_49 = ~(~n_585 | n_1073);
 assign sub_732_2_n_48 = ~(~n_661 | n_1105);
 assign sub_732_2_n_47 = ~(~n_697 & n_2397);
 assign sub_732_2_n_46 = ~(~n_1106 & n_1063);
 assign sub_732_2_n_45 = ~(~n_652 | n_2395);
 assign sub_732_2_n_44 = ~(~n_437 & n_2393);
 assign sub_732_2_n_43 = ~(~n_427 | n_2390);
 assign sub_732_2_n_42 = ~(~n_619 & n_1081);
 assign sub_732_2_n_41 = ~(~n_605 & n_1104);
 assign sub_732_2_n_40 = ~(~n_393 | n_2392);
 assign sub_732_2_n_39 = ~(~n_357 & n_2391);
 assign sub_732_2_n_38 = ~(~n_661 & n_1105);
 assign sub_732_2_n_37 = ~(~n_675 | n_2394);
 assign sub_732_2_n_36 = ~(~n_468 & n_2385);
 assign sub_732_2_n_35 = ~(~n_478 & n_2381);
 assign sub_732_2_n_34 = ~(n_468 & ~n_2385);
 assign sub_732_2_n_33 = ~({in1[0]} & ~{in2[1]});
 assign sub_732_2_n_32 = ~(~n_406 & n_1068);
 assign sub_732_2_n_31 = ~(n_406 & ~n_1068);
 assign sub_732_2_n_30 = ~(~n_634 & n_2396);
 assign sub_732_2_n_29 = ~(~n_530 & n_2398);
 assign sub_732_2_n_28 = ~(~n_530 | n_2398);
 assign sub_732_2_n_27 = ~(~n_1074 | n_457);
 assign sub_732_2_n_26 = ~(~n_1073 | n_585);
 assign sub_732_2_n_25 = ~(~n_560 & n_2384);
 assign sub_732_2_n_24 = ~(~n_1087 | n_549);
 assign sub_732_2_n_23 = ~(n_675 | ~n_2394);
 assign sub_732_2_n_22 = ~(~n_347 & n_2388);
 assign sub_732_2_n_21 = ~(~n_560 | n_2384);
 assign sub_732_2_n_20 = ~(~n_417 & n_2399);
 assign sub_732_2_n_19 = ~(~n_685 & n_2389);
 assign sub_732_2_n_18 = ~(~n_417 | n_2399);
 assign sub_732_2_n_17 = ~(n_1106 & ~n_1063);
 assign sub_732_2_n_16 = ~(~n_336 | n_2379);
 assign sub_732_2_n_15 = ~(~n_549 | n_1087);
 assign sub_732_2_n_14 = ~(~n_606 | n_2383);
 assign sub_732_2_n_13 = ~(~n_357 | n_2391);
 assign sub_732_2_n_12 = ~(~n_347 | n_2388);
 assign sub_732_2_n_11 = ~(~n_478 | n_2381);
 assign sub_732_2_n_10 = ~(~n_368 & n_2387);
 assign sub_732_2_n_9 = ~(~n_634 | n_2396);
 assign sub_732_2_n_8 = ~(~n_458 | n_2378);
 assign sub_732_2_n_7 = ~(~n_368 | n_2387);
 assign sub_732_2_n_6 = ~(~n_448 | n_2382);
 assign sub_732_2_n_5 = ~(~n_335 & n_1066);
 assign sub_732_2_n_4 = ~(~n_652 & n_2395);
 assign sub_732_2_n_3 = ~(n_697 & ~n_2397);
 assign sub_732_2_n_2 = ~(~n_437 | n_2393);
 assign sub_732_2_n_0 = (sub_732_2_n_62 | sub_732_2_n_43);
 assign n_2465 = ~(sub_751_2_n_71 ^ sub_751_2_n_199);
 assign sub_751_2_n_199 = ~(sub_751_2_n_52 & (sub_751_2_n_193 | sub_751_2_n_15));
 assign n_2473 = ~(sub_751_2_n_77 ^ sub_751_2_n_194);
 assign n_2466 = (sub_751_2_n_69 ^ sub_751_2_n_193);
 assign n_2467 = ~(sub_751_2_n_68 ^ sub_751_2_n_192);
 assign n_2469 = ~(sub_751_2_n_73 ^ sub_751_2_n_191);
 assign sub_751_2_n_194 = ~(sub_751_2_n_14 & (sub_751_2_n_183 | sub_751_2_n_6));
 assign sub_751_2_n_193 = ~(sub_751_2_n_112 | (sub_751_2_n_182 & sub_751_2_n_85));
 assign sub_751_2_n_192 = (~sub_751_2_n_10 | (sub_751_2_n_182 & sub_751_2_n_55));
 assign sub_751_2_n_191 = ~(sub_751_2_n_19 & (sub_751_2_n_178 | sub_751_2_n_5));
 assign n_2474 = (sub_751_2_n_96 ^ sub_751_2_n_183);
 assign n_2475 = (sub_751_2_n_99 ^ sub_751_2_n_180);
 assign n_2477 = ~(sub_751_2_n_95 ^ sub_751_2_n_179);
 assign n_2468 = ~(sub_751_2_n_67 ^ sub_751_2_n_182);
 assign n_2470 = (sub_751_2_n_64 ^ sub_751_2_n_178);
 assign n_2471 = ~(sub_751_2_n_75 ^ sub_751_2_n_173);
 assign n_2481 = (sub_751_2_n_88 ^ sub_751_2_n_172);
 assign n_2464 = (sub_751_2_n_140 & (sub_751_2_n_125 | n_3178));
 assign sub_751_2_n_180 = ~(sub_751_2_n_39 | (sub_751_2_n_168 & sub_751_2_n_56));
 assign sub_751_2_n_179 = ~(sub_751_2_n_41 & (sub_751_2_n_167 | sub_751_2_n_32));
 assign sub_751_2_n_183 = ~(sub_751_2_n_111 | (sub_751_2_n_168 & sub_751_2_n_106));
 assign sub_751_2_n_182 = ~(sub_751_2_n_130 & (n_3178 | sub_751_2_n_120));
 assign n_2476 = ~(sub_751_2_n_97 ^ sub_751_2_n_168);
 assign n_2472 = (sub_751_2_n_94 ^ n_3178);
 assign n_2479 = ~(sub_751_2_n_90 ^ sub_751_2_n_166);
 assign n_2478 = (sub_751_2_n_92 ^ sub_751_2_n_167);
 assign sub_751_2_n_173 = ~(sub_751_2_n_37 & (n_3178 | sub_751_2_n_11));
 assign sub_751_2_n_178 = (~sub_751_2_n_115 & (n_3178 | sub_751_2_n_105));
 assign sub_751_2_n_172 = ~(sub_751_2_n_38 | (sub_751_2_n_162 & sub_751_2_n_36));
 assign n_2482 = ~(sub_751_2_n_72 ^ sub_751_2_n_162);
 assign n_2483 = (sub_751_2_n_87 ^ sub_751_2_n_161);
 assign n_2485 = (sub_751_2_n_98 ^ sub_751_2_n_160);
 assign sub_751_2_n_168 = ~(sub_751_2_n_131 & (sub_751_2_n_156 | sub_751_2_n_118));
 assign sub_751_2_n_167 = (~sub_751_2_n_113 & (sub_751_2_n_156 | sub_751_2_n_109));
 assign sub_751_2_n_166 = ~(sub_751_2_n_34 & (sub_751_2_n_156 | sub_751_2_n_13));
 assign n_2480 = (sub_751_2_n_89 ^ sub_751_2_n_156);
 assign sub_751_2_n_162 = ~(sub_751_2_n_117 & (sub_751_2_n_155 | sub_751_2_n_110));
 assign sub_751_2_n_161 = (~sub_751_2_n_2 & (sub_751_2_n_155 | sub_751_2_n_42));
 assign sub_751_2_n_160 = ~(sub_751_2_n_46 | (sub_751_2_n_154 & sub_751_2_n_40));
 assign n_2484 = (sub_751_2_n_93 ^ sub_751_2_n_155);
 assign n_2486 = ~(sub_751_2_n_66 ^ sub_751_2_n_154);
 assign n_2487 = (sub_751_2_n_91 ^ sub_751_2_n_153);
 assign sub_751_2_n_156 = ~(sub_751_2_n_138 | (sub_751_2_n_150 & (sub_751_2_n_123 & sub_751_2_n_122)));
 assign sub_751_2_n_155 = ~(sub_751_2_n_132 | (sub_751_2_n_150 & sub_751_2_n_122));
 assign sub_751_2_n_154 = (~sub_751_2_n_116 | (sub_751_2_n_150 & sub_751_2_n_104));
 assign sub_751_2_n_153 = ~(sub_751_2_n_49 | (sub_751_2_n_150 & sub_751_2_n_47));
 assign n_2488 = ~(sub_751_2_n_70 ^ sub_751_2_n_150);
 assign n_2489 = ~(sub_751_2_n_62 ^ sub_751_2_n_149);
 assign sub_751_2_n_150 = ~(sub_751_2_n_145 & (sub_751_2_n_29 & sub_751_2_n_129));
 assign sub_751_2_n_149 = ~(sub_751_2_n_9 & (sub_751_2_n_146 | sub_751_2_n_20));
 assign n_2490 = (sub_751_2_n_76 ^ sub_751_2_n_146);
 assign n_2491 = ~(sub_751_2_n_74 ^ sub_751_2_n_144);
 assign sub_751_2_n_146 = ~(sub_751_2_n_114 | (sub_751_2_n_142 & sub_751_2_n_82));
 assign sub_751_2_n_145 = ~(sub_751_2_n_142 & (sub_751_2_n_80 & sub_751_2_n_82));
 assign sub_751_2_n_144 = (~sub_751_2_n_4 | (sub_751_2_n_142 & sub_751_2_n_7));
 assign n_2492 = (sub_751_2_n_63 ^ sub_751_2_n_142);
 assign sub_751_2_n_142 = ~(sub_751_2_n_30 & (sub_751_2_n_27 | (sub_751_2_n_135 & sub_751_2_n_17)));
 assign n_2493 = (sub_751_2_n_65 ^ sub_751_2_n_139);
 assign sub_751_2_n_140 = (sub_751_2_n_31 & (sub_751_2_n_128 & (sub_751_2_n_130 | sub_751_2_n_119)));
 assign sub_751_2_n_139 = (sub_751_2_n_17 & ~(sub_751_2_n_134 & sub_751_2_n_33));
 assign sub_751_2_n_138 = (sub_751_2_n_26 | (sub_751_2_n_127 | (sub_751_2_n_132 & sub_751_2_n_123)));
 assign sub_751_2_n_137 = ~(sub_751_2_n_59 & (sub_751_2_n_126 & (sub_751_2_n_131 | sub_751_2_n_121)));
 assign n_2494 = (sub_751_2_n_134 ^ sub_751_2_n_100);
 assign sub_751_2_n_135 = ~(sub_751_2_n_134 & sub_751_2_n_33);
 assign sub_751_2_n_134 = ((n_382 & n_497) | (n_2463 & (n_382 ^ n_497)));
 assign n_2495 = (n_2463 ^ (n_382 ^ n_497));
 assign sub_751_2_n_132 = ~(sub_751_2_n_101 & (sub_751_2_n_25 & (sub_751_2_n_116 | sub_751_2_n_107)));
 assign sub_751_2_n_131 = ~(sub_751_2_n_79 | (sub_751_2_n_60 | (sub_751_2_n_113 & sub_751_2_n_83)));
 assign sub_751_2_n_130 = ~(sub_751_2_n_103 | (sub_751_2_n_22 | (sub_751_2_n_115 & sub_751_2_n_84)));
 assign sub_751_2_n_129 = ~((~sub_751_2_n_9 & ~sub_751_2_n_51) | (sub_751_2_n_114 & sub_751_2_n_80));
 assign sub_751_2_n_128 = ~((~sub_751_2_n_52 & ~sub_751_2_n_54) | (sub_751_2_n_112 & sub_751_2_n_86));
 assign sub_751_2_n_127 = ~(sub_751_2_n_102 & (sub_751_2_n_117 | sub_751_2_n_81));
 assign sub_751_2_n_126 = ~((~sub_751_2_n_14 & ~sub_751_2_n_3) | (sub_751_2_n_111 & sub_751_2_n_108));
 assign sub_751_2_n_125 = (sub_751_2_n_120 | sub_751_2_n_119);
 assign sub_751_2_n_124 = (sub_751_2_n_118 | sub_751_2_n_121);
 assign sub_751_2_n_123 = ~(sub_751_2_n_110 | sub_751_2_n_81);
 assign sub_751_2_n_122 = ~(sub_751_2_n_107 | ~sub_751_2_n_104);
 assign sub_751_2_n_121 = ~(sub_751_2_n_106 & sub_751_2_n_108);
 assign sub_751_2_n_120 = ~(~sub_751_2_n_105 & sub_751_2_n_84);
 assign sub_751_2_n_119 = ~(sub_751_2_n_85 & sub_751_2_n_86);
 assign sub_751_2_n_118 = ~(~sub_751_2_n_109 & sub_751_2_n_83);
 assign sub_751_2_n_117 = ~(sub_751_2_n_21 | (sub_751_2_n_2 & sub_751_2_n_35));
 assign sub_751_2_n_116 = ~(sub_751_2_n_57 | (sub_751_2_n_49 & sub_751_2_n_44));
 assign sub_751_2_n_115 = ~(sub_751_2_n_58 & (sub_751_2_n_37 | sub_751_2_n_48));
 assign sub_751_2_n_114 = ~(sub_751_2_n_24 & (sub_751_2_n_4 | sub_751_2_n_53));
 assign sub_751_2_n_113 = ~(sub_751_2_n_28 & (sub_751_2_n_34 | sub_751_2_n_12));
 assign sub_751_2_n_112 = ~(sub_751_2_n_23 & (sub_751_2_n_10 | sub_751_2_n_16));
 assign sub_751_2_n_111 = (~sub_751_2_n_61 | (sub_751_2_n_39 & sub_751_2_n_45));
 assign sub_751_2_n_103 = ~(sub_751_2_n_19 | sub_751_2_n_43);
 assign sub_751_2_n_102 = ~(sub_751_2_n_38 & sub_751_2_n_8);
 assign sub_751_2_n_101 = ~(sub_751_2_n_46 & sub_751_2_n_18);
 assign sub_751_2_n_110 = ~(~sub_751_2_n_42 & sub_751_2_n_35);
 assign sub_751_2_n_100 = (sub_751_2_n_17 & sub_751_2_n_33);
 assign sub_751_2_n_99 = ~(sub_751_2_n_61 & sub_751_2_n_45);
 assign sub_751_2_n_98 = ~(sub_751_2_n_25 & sub_751_2_n_18);
 assign sub_751_2_n_97 = ~(sub_751_2_n_56 & ~sub_751_2_n_39);
 assign sub_751_2_n_109 = (sub_751_2_n_13 | sub_751_2_n_12);
 assign sub_751_2_n_108 = ~(sub_751_2_n_6 | sub_751_2_n_3);
 assign sub_751_2_n_96 = ~(sub_751_2_n_14 & ~sub_751_2_n_6);
 assign sub_751_2_n_95 = ~(sub_751_2_n_50 & ~sub_751_2_n_60);
 assign sub_751_2_n_94 = ~(sub_751_2_n_37 & ~sub_751_2_n_11);
 assign sub_751_2_n_93 = (sub_751_2_n_2 | sub_751_2_n_42);
 assign sub_751_2_n_92 = ~(~sub_751_2_n_32 & sub_751_2_n_41);
 assign sub_751_2_n_91 = ~(sub_751_2_n_44 & ~sub_751_2_n_57);
 assign sub_751_2_n_107 = ~(sub_751_2_n_40 & sub_751_2_n_18);
 assign sub_751_2_n_90 = ~(sub_751_2_n_28 & ~sub_751_2_n_12);
 assign sub_751_2_n_106 = (sub_751_2_n_56 & sub_751_2_n_45);
 assign sub_751_2_n_105 = (sub_751_2_n_11 | sub_751_2_n_48);
 assign sub_751_2_n_89 = ~(sub_751_2_n_34 & ~sub_751_2_n_13);
 assign sub_751_2_n_88 = ~(sub_751_2_n_8 & ~sub_751_2_n_26);
 assign sub_751_2_n_104 = (sub_751_2_n_47 & sub_751_2_n_44);
 assign sub_751_2_n_87 = ~(sub_751_2_n_35 & ~sub_751_2_n_21);
 assign sub_751_2_n_79 = ~(sub_751_2_n_41 | ~sub_751_2_n_50);
 assign n_2496 = ~(sub_751_2_n_1 & (~{in2[0]} | {in1[0]}));
 assign sub_751_2_n_77 = ~(sub_751_2_n_59 & ~sub_751_2_n_3);
 assign sub_751_2_n_76 = ~(~sub_751_2_n_20 & sub_751_2_n_9);
 assign sub_751_2_n_75 = ~(sub_751_2_n_58 & ~sub_751_2_n_48);
 assign sub_751_2_n_74 = ~(sub_751_2_n_24 & ~sub_751_2_n_53);
 assign sub_751_2_n_73 = (sub_751_2_n_22 | sub_751_2_n_43);
 assign sub_751_2_n_86 = ~(sub_751_2_n_15 | sub_751_2_n_54);
 assign sub_751_2_n_72 = ~(sub_751_2_n_36 & ~sub_751_2_n_38);
 assign sub_751_2_n_85 = ~(sub_751_2_n_16 | ~sub_751_2_n_55);
 assign sub_751_2_n_71 = ~(sub_751_2_n_31 & ~sub_751_2_n_54);
 assign sub_751_2_n_84 = ~(sub_751_2_n_5 | sub_751_2_n_43);
 assign sub_751_2_n_70 = ~(sub_751_2_n_47 & ~sub_751_2_n_49);
 assign sub_751_2_n_69 = ~(sub_751_2_n_52 & ~sub_751_2_n_15);
 assign sub_751_2_n_68 = ~(sub_751_2_n_23 & ~sub_751_2_n_16);
 assign sub_751_2_n_83 = ~(sub_751_2_n_32 | ~sub_751_2_n_50);
 assign sub_751_2_n_67 = ~(sub_751_2_n_10 & sub_751_2_n_55);
 assign sub_751_2_n_66 = ~(sub_751_2_n_40 & ~sub_751_2_n_46);
 assign sub_751_2_n_82 = ~(sub_751_2_n_53 | ~sub_751_2_n_7);
 assign sub_751_2_n_65 = ~(sub_751_2_n_30 & ~sub_751_2_n_27);
 assign sub_751_2_n_81 = ~(sub_751_2_n_36 & sub_751_2_n_8);
 assign sub_751_2_n_64 = ~(sub_751_2_n_19 & ~sub_751_2_n_5);
 assign sub_751_2_n_63 = (sub_751_2_n_4 & sub_751_2_n_7);
 assign sub_751_2_n_62 = ~(sub_751_2_n_29 & ~sub_751_2_n_51);
 assign sub_751_2_n_80 = ~(sub_751_2_n_20 | sub_751_2_n_51);
 assign sub_751_2_n_61 = ~(~n_595 & n_2443);
 assign sub_751_2_n_60 = ~(~n_2445 | n_447);
 assign sub_751_2_n_59 = ~(~n_457 & n_2441);
 assign sub_751_2_n_58 = ~(~n_539 & n_2439);
 assign sub_751_2_n_57 = ~(~n_2455 | n_392);
 assign sub_751_2_n_56 = ~(n_477 & ~n_2444);
 assign sub_751_2_n_55 = ~(~n_2436 & n_619);
 assign sub_751_2_n_54 = ~(~n_498 | n_2433);
 assign sub_751_2_n_53 = ~(~n_633 | n_2459);
 assign sub_751_2_n_52 = ~(~n_406 & n_2434);
 assign sub_751_2_n_51 = ~(~n_674 | n_2457);
 assign sub_751_2_n_50 = ~(n_447 & ~n_2445);
 assign sub_751_2_n_49 = ~(~n_2456 | n_436);
 assign sub_751_2_n_48 = ~(~n_539 | n_2439);
 assign sub_751_2_n_47 = ~(n_436 & ~n_2456);
 assign sub_751_2_n_46 = ~(~n_2454 | n_356);
 assign sub_751_2_n_45 = ~(n_595 & ~n_2443);
 assign sub_751_2_n_44 = ~(~n_2455 & n_392);
 assign sub_751_2_n_43 = ~(~n_549 | n_2437);
 assign sub_751_2_n_42 = ~(~n_684 | n_2452);
 assign sub_751_2_n_41 = ~(~n_605 & n_2446);
 assign sub_751_2_n_40 = ~(~n_2454 & n_356);
 assign sub_751_2_n_39 = ~(~n_2444 | n_477);
 assign sub_751_2_n_38 = ~(~n_2450 | n_367);
 assign sub_751_2_n_37 = ~(~n_1106 & n_2440);
 assign sub_751_2_n_36 = ~(~n_2450 & n_367);
 assign sub_751_2_n_35 = ~(~n_2451 & n_346);
 assign sub_751_2_n_34 = ~(~n_467 & n_2448);
 assign sub_751_2_n_33 = ~(~n_2462 & n_416);
 assign sub_751_2_n_32 = ~(~n_605 | n_2446);
 assign sub_751_2_n_31 = ~(~n_498 & n_2433);
 assign sub_751_2_n_30 = ~(~n_529 & n_2461);
 assign sub_751_2_n_29 = ~(~n_674 & n_2457);
 assign sub_751_2_n_28 = ~(~n_559 & n_2447);
 assign sub_751_2_n_27 = ~(~n_529 | n_2461);
 assign sub_751_2_n_26 = ~(~n_2449 | n_518);
 assign sub_751_2_n_25 = ~(~n_426 & n_2453);
 assign sub_751_2_n_24 = ~(~n_633 & n_2459);
 assign sub_751_2_n_23 = ~(~n_585 & n_2435);
 assign sub_751_2_n_22 = ~(~n_2437 | n_549);
 assign sub_751_2_n_21 = ~(~n_2451 | n_346);
 assign sub_751_2_n_20 = ~(~n_651 | n_2458);
 assign sub_751_2_n_19 = ~(~n_661 & n_2438);
 assign sub_751_2_n_18 = ~(~n_2453 & n_426);
 assign sub_751_2_n_17 = ~(~n_416 & n_2462);
 assign sub_751_2_n_16 = ~(~n_585 | n_2435);
 assign sub_751_2_n_15 = ~(~n_406 | n_2434);
 assign sub_751_2_n_14 = ~(~n_335 & n_2442);
 assign sub_751_2_n_13 = ~(~n_467 | n_2448);
 assign sub_751_2_n_12 = ~(~n_559 | n_2447);
 assign sub_751_2_n_11 = ~(~n_1106 | n_2440);
 assign sub_751_2_n_10 = ~(~n_619 & n_2436);
 assign sub_751_2_n_9 = ~(~n_651 & n_2458);
 assign sub_751_2_n_8 = ~(~n_2449 & n_518);
 assign sub_751_2_n_7 = ~(n_696 & ~n_2460);
 assign sub_751_2_n_6 = ~(~n_335 | n_2442);
 assign sub_751_2_n_5 = ~(~n_661 | n_2438);
 assign sub_751_2_n_4 = ~(~n_696 & n_2460);
 assign sub_751_2_n_3 = ~(~n_457 | n_2441);
 assign sub_751_2_n_2 = ~(~n_2452 | n_684);
 assign sub_751_2_n_1 = ~({in1[0]} & ~{in2[0]});
 assign sub_751_2_n_0 = ~n_383;
 assign n_268 = ~clr;
 assign n_3042 = ((n_726 & ~n_2554) | (n_725 & n_2554));
 assign n_3043 = ((n_1511 & ~n_1504) | (n_3042 & n_1504));
 assign n_3044 = ((n_712 & ~n_1521) | (n_713 & n_1521));
 assign n_3045 = ((n_1547 & ~n_1540) | (n_749 & n_1540));
 assign n_3038 = ((n_577 & ~n_1540) | (n_578 & n_1540));
 assign n_3047 = ((n_1546 & ~n_1540) | (n_734 & n_1540));
 assign n_3048 = ((n_1569 & ~n_1561) | (n_3245 & n_1561));
 assign n_3049 = ((n_580 & ~n_1584) | (n_581 & n_1584));
 assign n_3050 = ((n_582 & ~n_780) | (n_584 & n_780));
 assign n_3051 = ((n_630 & ~n_1636) | (n_632 & n_1636));
 assign n_3052 = ((n_1649 & ~n_1636) | (n_3050 & n_1636));
 assign n_3053 = ((n_3279 & ~n_2677) | (n_1666 & n_2677));
 assign n_3054 = ((n_1652 & ~n_2677) | (n_1667 & n_2677));
 assign n_3055 = ((n_787 & ~n_2717) | (n_789 & n_2717));
 assign n_3056 = ((n_785 & ~n_1729) | (n_786 & n_1729));
 assign n_3057 = ((n_490 & ~n_1729) | (n_492 & n_1729));
 assign n_3058 = ((n_403 & ~n_1764) | (n_405 & n_1764));
 assign n_3059 = ((n_650 & ~n_1801) | (n_671 & n_1801));
 assign n_3060 = ((n_2089 & ~n_2065) | (n_926 & n_2065));
 assign n_3061 = ((n_377 & ~n_2065) | (n_345 & n_2065));
 assign n_3062 = ((n_2141 & ~n_2116) | (n_3061 & n_2116));
 assign n_3063 = ((n_446 & ~n_2116) | (n_720 & n_2116));
 assign n_3064 = ((n_570 & ~n_2169) | (n_573 & n_2169));
 assign n_3065 = ((n_960 & ~n_2169) | (n_961 & n_2169));
 assign n_3066 = ((n_1003 & ~n_2169) | (n_1007 & n_2169));
 assign n_3067 = ((n_957 & ~n_2169) | (n_950 & n_2169));
 assign n_3068 = ((n_2251 & ~n_2224) | (n_3064 & n_2224));
 assign n_3070 = ~({in1[1]} | (n_3069 | ~n_3117));
 assign n_3069 = ~(n_3106 & (n_3717 & n_3716));
 assign n_3071 = ~(sub_219_2_n_4 ^ (n_3221 ^ {in1[1]}));
 assign n_3072 = ~({in1[8]} | ({in1[9]} | ({in1[10]} | {in1[11]})));
 assign n_3080 = ~({in1[10]} | {in1[11]});
 assign n_3083 = ~({in1[8]} | {in1[9]});
 assign n_3092 = ~({in1[28]} | {in1[29]});
 assign n_3095 = ~({in1[26]} | {in1[27]});
 assign n_3099 = ~({in1[24]} | {in1[25]});
 assign n_3102 = ~({in1[22]} | {in1[23]});
 assign n_3105 = ~({in1[20]} | {in1[21]});
 assign n_3106 = ~({in1[2]} | {in1[3]});
 assign n_3109 = ~({in1[12]} | {in1[13]});
 assign n_3113 = ~({in1[6]} | {in1[7]});
 assign n_3117 = ~({in1[18]} | {in1[19]});
 assign n_3118 = ~({in1[26]} | ({in1[27]} | ({in1[28]} | {in1[29]})));
 assign n_3119 = ~({in1[20]} | ({in1[21]} | ({in1[22]} | {in1[23]})));
 assign n_3121 = ~(n_486 | (n_604 | (n_344 | n_466)));
 assign n_3122 = ~(n_614 | n_456);
 assign n_3123 = ~(n_376 | (n_527 | (n_476 | n_568)));
 assign n_3124 = ~(n_693 | n_355);
 assign n_3125 = ~(n_445 | (n_401 | (n_365 | n_435)));
 assign n_3126 = ~(n_415 | n_507);
 assign n_3127 = ~(n_670 | (n_558 | (n_628 | n_594)));
 assign n_3128 = ~(n_1115 | n_548);
 assign n_3129 = ~(n_692 | (n_354 | (n_375 | n_526)));
 assign n_3131 = ~(n_475 | n_567);
 assign n_3134 = ~(n_485 | (n_603 | (n_343 | n_465)));
 assign n_3136 = ~(n_627 | (n_593 | (n_414 | n_506)));
 assign n_3137 = ~(n_547 | n_669);
 assign n_3138 = ~(n_484 | n_602);
 assign n_3139 = ~(n_474 | (n_566 | (n_612 | n_454)));
 assign n_3140 = ~(n_546 | n_668);
 assign n_3141 = ~(n_626 | (n_592 | (n_413 | n_505)));
 assign n_3142 = ~(n_625 | n_504);
 assign n_3143 = ~(n_1112 | (n_545 | (n_667 | n_555)));
 assign n_3144 = ~(n_483 | (n_601 | (n_341 | n_463)));
 assign n_3145 = ~(n_611 | n_453);
 assign n_3146 = ~(n_1111 | n_554);
 assign n_3147 = ~(n_624 | (n_590 | (n_411 | n_503)));
 assign n_3148 = ~(n_340 | n_462);
 assign n_3149 = ~(n_665 | n_553);
 assign n_3150 = ~(n_623 | (n_589 | (n_410 | n_502)));
 assign n_3152 = ~(n_1110 | n_543);
 assign n_3153 = ~(n_664 | n_552);
 assign n_3154 = (n_622 | (n_588 | (n_409 | n_501)));
 assign n_3159 = ~(n_3105 & (n_3102 & n_3099));
 assign n_3161 = ~(n_3083 & (n_3080 & n_3109));
 assign n_3164 = ~(n_3119 & (n_3099 & (n_3118 & n_3718)));
 assign n_3165 = ~(n_3125 & (n_3124 & (n_3123 & n_3122)));
 assign n_3166 = ~(n_3121 & (n_3128 & (n_3127 & n_3126)));
 assign n_3167 = ~(~n_3136 | (n_1114 | n_557));
 assign n_3169 = ~(n_3201 & (~sub_333_2_n_0 & ~n_3544));
 assign n_3170 = ~(n_3167 & (n_3137 & (n_3134 & n_3131)));
 assign n_3171 = ~(sub_466_2_n_110 & (~n_804 & ~sub_466_2_n_96));
 assign n_3172 = ~(n_613 | (n_455 | n_3170));
 assign n_3173 = ~(~n_423 | n_3272);
 assign n_3174 = ~(~n_691 & n_3268);
 assign n_3175 = ~(sub_409_2_n_89 & (~sub_409_2_n_43 & ~sub_409_2_n_78));
 assign n_3176 = ~(~n_444 & n_3249);
 assign n_3177 = ~(sub_675_2_n_154 & (~sub_675_2_n_52 & ~sub_675_2_n_138));
 assign n_3178 = (~sub_751_2_n_137 & (sub_751_2_n_156 | sub_751_2_n_124));
 assign n_3179 = ~(~sub_675_2_n_135 & sub_675_2_n_169);
 assign n_3180 = ~(~n_363 & n_3278);
 assign n_3181 = ~(~sub_675_2_n_148 & n_3179);
 assign n_3182 = ~(~n_691 & n_3280);
 assign n_3183 = ~(~{in1[2]} & n_3220);
 assign n_3185 = ~(sub_371_2_n_81 & (~sub_371_2_n_45 & ~sub_371_2_n_70));
 assign n_3188 = ~(~n_424 | n_1607);
 assign n_3189 = ~(sub_447_2_n_16 | (~sub_447_2_n_94 & sub_447_2_n_19));
 assign n_3190 = ~(~n_640 | n_3306);
 assign n_3192 = (n_644 ^ sub_276_2_n_27);
 assign n_3193 = (n_645 ^ sub_314_2_n_39);
 assign n_3194 = ~(n_538 & ~n_1537);
 assign n_3197 = ~(sub_257_2_n_44 & (n_3113 & ~sub_257_2_n_35));
 assign n_3199 = ~(sub_314_2_n_35 & (~sub_314_2_n_42 | sub_314_2_n_44));
 assign n_3200 = ~(n_705 | ~n_3723);
 assign n_3201 = ~(n_745 & (n_740 & n_739));
 assign n_3202 = ~(sub_352_2_n_78 & (sub_352_2_n_4 & ~sub_352_2_n_61));
 assign n_3036 = ~(~n_659 & n_3246);
 assign n_3204 = ~(sub_390_2_n_8 | (~sub_390_2_n_38 & sub_390_2_n_1));
 assign n_3205 = ~(~n_424 & n_1607);
 assign n_3207 = ~(~n_3293 & n_536);
 assign n_3208 = ~(~n_681 & n_3291);
 assign n_3209 = ~(n_640 | ~n_3306);
 assign n_3210 = (sub_485_2_n_58 & ~(sub_485_2_n_9 & sub_485_2_n_104));
 assign n_3211 = ~(~n_3317 & n_690);
 assign n_3212 = ~(sub_561_2_n_104 | (sub_561_2_n_83 & sub_561_2_n_139));
 assign n_3213 = ~(n_386 | ~n_3425);
 assign n_3214 = ~(~n_3513 & n_531);
 assign n_3216 = ~n_3215;
 assign n_3215 = ~({in2[31]} & (~{in1[0]} | n_1441));
 assign n_3217 = (~n_2502 | (n_1445 & n_2503));
 assign n_3218 = ((n_3536 & n_2503) | (n_1444 & {in2[30]}));
 assign n_3219 = ((n_1450 & n_2511) | (n_3217 & n_1449));
 assign n_3220 = ((n_1451 & n_2511) | (n_3218 & n_1449));
 assign n_3221 = (~n_3222 | (n_1449 & {in2[29]}));
 assign n_3222 = (~n_2511 | (sub_200_2_n_2 & sub_200_2_n_6));
 assign n_3223 = ((n_1457 & n_2521) | (n_3219 & n_2519));
 assign n_3224 = (~n_2516 | (n_1460 & n_2520));
 assign n_3225 = (~n_2536 | (n_1465 & {in2[27]}));
 assign n_3226 = ((n_1467 & n_2532) | (n_3228 & n_1465));
 assign n_3227 = ((n_1492 & n_2554) | (n_3236 & n_2553));
 assign n_3228 = ((n_1458 & n_2521) | (n_3220 & n_2519));
 assign n_3229 = ((n_3071 & n_2520) | (n_3221 & n_2522));
 assign n_3230 = ((n_1466 & n_2532) | (n_3223 & n_1465));
 assign n_3231 = ((n_1469 & n_2532) | (n_3224 & n_1465));
 assign n_3232 = ((n_1477 & n_2542) | (n_711 & n_1476));
 assign n_3233 = ((n_721 & n_2542) | (n_724 & n_1476));
 assign n_3234 = ((n_647 & n_2542) | (n_649 & n_1476));
 assign n_3235 = ((n_694 & n_2542) | (n_648 & n_1476));
 assign n_3236 = ((n_718 & n_2542) | (n_646 & n_1476));
 assign n_3237 = ((n_617 & n_2542) | (n_1476 & n_643));
 assign n_3238 = ((n_1490 & n_2554) | (n_3232 & n_2553));
 assign n_3239 = ((n_1491 & n_2554) | (n_3235 & n_2553));
 assign n_3240 = ((n_1494 & n_2554) | (n_3234 & n_2553));
 assign n_3241 = ((n_1508 & n_2567) | (n_1500 & n_1504));
 assign n_3242 = ((n_2567 & n_488) | (n_1504 & n_489));
 assign n_3243 = ((n_1544 & n_2590) | (n_750 & n_1540));
 assign n_3244 = ((n_2590 & n_1541) | (n_727 & n_1540));
 assign n_3245 = ((n_1548 & n_2590) | (n_747 & n_1540));
 assign n_3246 = ((n_1545 & n_2590) | (n_742 & n_1540));
 assign n_3247 = ((n_1542 & n_2590) | (n_743 & n_1540));
 assign n_3248 = (~n_2600 | (n_737 & n_1540));
 assign n_3249 = ((n_1543 & n_2590) | (n_738 & n_1540));
 assign n_3250 = ((n_2607 & n_1562) | (n_3244 & n_2606));
 assign n_3251 = ((n_2607 & n_1563) | (n_3247 & n_2606));
 assign n_3252 = ((n_1564 & n_2607) | (n_3249 & n_2606));
 assign n_3253 = ((n_1567 & n_2607) | (n_3047 & n_1561));
 assign n_3254 = ((n_2623 & n_1585) | (n_3250 & n_2624));
 assign n_3255 = ((n_1588 & n_2623) | (n_1576 & n_2624));
 assign n_3256 = ((n_1591 & n_2623) | (n_1579 & n_1584));
 assign n_3257 = ((n_2623 & n_1592) | (n_3048 & n_1584));
 assign n_3258 = ((n_2623 & n_1593) | (n_3726 & n_1584));
 assign n_3259 = ((n_1594 & n_2623) | (n_3727 & n_1584));
 assign n_3260 = ((n_2623 & n_1586) | (n_3251 & n_2624));
 assign n_3261 = ((n_1590 & n_2623) | (n_3253 & n_1584));
 assign n_3262 = ((n_2637 & n_1610) | (n_774 & n_780));
 assign n_3263 = ((n_2637 & n_1613) | (n_763 & n_780));
 assign n_3264 = ((n_757 & n_2637) | (n_778 & n_780));
 assign n_3265 = ((n_756 & n_2637) | (n_779 & n_780));
 assign n_3266 = ((n_770 & n_2637) | (n_773 & n_780));
 assign n_3267 = ((n_2637 & n_755) | (n_777 & n_780));
 assign n_3268 = ((n_2637 & n_1611) | (n_752 & n_780));
 assign n_3269 = ((n_2637 & n_1612) | (n_767 & n_780));
 assign n_3270 = ((n_2637 & n_760) | (n_761 & n_780));
 assign n_3271 = ((n_753 & n_2637) | (n_776 & n_780));
 assign n_3272 = ((n_754 & n_2637) | (n_775 & n_780));
 assign n_3273 = ((n_758 & n_2637) | (n_759 & n_780));
 assign n_3274 = ((n_1645 & n_2658) | (n_3267 & n_1636));
 assign n_3275 = ((n_2658 & n_1640) | (n_3263 & n_2657));
 assign n_3276 = ((n_2658 & n_1643) | (n_3264 & n_2657));
 assign n_3277 = ((n_1644 & n_2658) | (n_3265 & n_1636));
 assign n_3278 = ((n_2658 & n_1641) | (n_3266 & n_2657));
 assign n_3279 = ((n_2658 & n_1637) | (n_3262 & n_2657));
 assign n_3280 = ((n_2658 & n_1639) | (n_3269 & n_2657));
 assign n_3281 = ((n_2658 & n_1642) | (n_3270 & n_2657));
 assign n_3282 = ((n_1647 & n_2658) | (n_3271 & n_1636));
 assign n_3283 = ((n_1648 & n_2658) | (n_3272 & n_1636));
 assign n_3284 = ((n_1646 & n_2658) | (n_3273 & n_1636));
 assign n_3285 = ((n_2677 & n_1670) | (n_3278 & n_1665));
 assign n_3286 = ((n_2677 & n_1669) | (n_3275 & n_1665));
 assign n_3287 = ((n_1672 & n_2677) | (n_3276 & n_1665));
 assign n_3288 = ((n_2677 & n_1679) | (n_3051 & n_1665));
 assign n_3289 = ((n_2677 & n_1671) | (n_3281 & n_1665));
 assign n_3290 = ((n_2677 & n_1668) | (n_3280 & n_1665));
 assign n_3291 = ((n_1674 & n_2677) | (n_3274 & n_1665));
 assign n_3292 = ((n_1676 & n_2677) | (n_3282 & n_1665));
 assign n_3293 = ((n_2677 & n_1678) | (n_3052 & n_1665));
 assign n_3294 = ((n_2696 & n_1704) | (n_1688 & n_1696));
 assign n_3295 = ((n_2696 & n_1700) | (n_3286 & n_1696));
 assign n_3296 = ((n_2696 & n_1703) | (n_3287 & n_1696));
 assign n_3297 = ((n_1710 & n_2696) | (n_3288 & n_1696));
 assign n_3298 = ((n_2696 & n_1697) | (n_3053 & n_1696));
 assign n_3299 = ((n_2696 & n_1701) | (n_3285 & n_1696));
 assign n_3300 = ((n_2696 & n_1702) | (n_3289 & n_1696));
 assign n_3301 = ((n_1706 & n_2696) | (n_1690 & n_1696));
 assign n_3302 = ((n_2696 & n_1698) | (n_3054 & n_1696));
 assign n_3303 = ((n_2696 & n_1699) | (n_3290 & n_1696));
 assign n_3304 = ((n_1705 & n_2696) | (n_3291 & n_1696));
 assign n_3305 = ((n_1707 & n_2696) | (n_3292 & n_1696));
 assign n_3306 = ((n_1708 & n_2696) | (n_1692 & n_1696));
 assign n_3307 = ((n_2719 & n_1737) | (n_821 & n_2717));
 assign n_3308 = ((n_2719 & n_1733) | (n_832 & n_2717));
 assign n_3309 = ((n_1736 & n_2719) | (n_820 & n_2717));
 assign n_3312 = ((n_1734 & n_2719) | (n_828 & n_2717));
 assign n_3314 = ((n_2719 & n_1739) | (n_805 & n_2717));
 assign n_3316 = ((n_2719 & n_1732) | (n_799 & n_2717));
 assign n_3317 = ((n_2719 & n_1735) | (n_783 & n_2717));
 assign n_3318 = ((n_1740 & n_2719) | (n_794 & n_2717));
 assign n_3319 = ((n_1741 & n_2719) | (n_827 & n_2717));
 assign n_3320 = ((n_2719 & n_1738) | (n_795 & n_2717));
 assign n_3321 = ((n_1768 & n_2747) | (n_3308 & n_2748));
 assign n_3322 = ((n_2747 & n_1778) | (n_3728 & n_1764));
 assign n_3323 = ((n_1780 & n_2747) | (n_3056 & n_1764));
 assign n_3324 = ((n_2747 & n_1769) | (n_3312 & n_2748));
 assign n_3325 = ((n_2747 & n_1777) | (n_3730 & n_1764));
 assign n_3326 = ((n_2747 & n_1774) | (n_3314 & n_1764));
 assign n_3327 = ((n_2749 & n_1766) | (n_3731 & n_2748));
 assign n_3328 = ((n_2749 & n_1767) | (n_3316 & n_2748));
 assign n_3329 = ((n_1775 & n_2747) | (n_3318 & n_1764));
 assign n_3330 = ((n_2747 & n_1776) | (n_3319 & n_1764));
 assign n_3331 = ((n_2781 & n_1817) | (n_3323 & n_1801));
 assign n_3332 = ((n_2781 & n_1806) | (n_3324 & n_1801));
 assign n_3333 = ((n_2781 & n_1802) | (n_1783 & n_1801));
 assign n_3337 = ((n_2781 & n_1803) | (n_3327 & n_1801));
 assign n_3338 = ((n_2781 & n_1804) | (n_3328 & n_1801));
 assign n_3339 = ((n_2781 & n_1807) | (n_1788 & n_1801));
 assign n_3341 = ((n_2781 & n_1813) | (n_3330 & n_1801));
 assign n_3343 = ((n_2805 & n_1841) | (n_849 & n_3699));
 assign n_3344 = ((n_2805 & n_1844) | (n_846 & n_3699));
 assign n_3345 = ((n_2805 & n_1847) | (n_836 & n_3699));
 assign n_3346 = ((n_2805 & n_1854) | (n_845 & n_3699));
 assign n_3347 = ((n_2805 & n_1848) | (n_835 & n_3699));
 assign n_3348 = ((n_2805 & n_1855) | (n_838 & n_3699));
 assign n_3349 = ((n_2805 & n_1856) | (n_852 & n_3699));
 assign n_3350 = ((n_2805 & n_1845) | (n_850 & n_3699));
 assign n_3351 = ((n_2805 & n_1849) | (n_833 & n_3699));
 assign n_3352 = ((n_2805 & n_1857) | (n_841 & n_3699));
 assign n_3353 = ((n_2805 & n_1858) | (n_842 & n_3699));
 assign n_3354 = ((n_2805 & n_1850) | (n_834 & n_3699));
 assign n_3355 = ((n_2805 & n_839) | (n_843 & n_3699));
 assign n_3356 = ((n_2805 & n_1842) | (n_851 & n_3699));
 assign n_3357 = ((n_2805 & n_1843) | (n_853 & n_3699));
 assign n_3358 = ((n_2805 & n_575) | (n_3699 & n_629));
 assign n_3359 = ((n_2805 & n_1846) | (n_848 & n_3699));
 assign n_3360 = ((n_2805 & n_1851) | (n_837 & n_3699));
 assign n_3361 = ((n_2805 & n_1852) | (n_847 & n_3699));
 assign n_3362 = ((n_2805 & n_1853) | (n_844 & n_3699));
 assign n_3363 = ((n_2833 & n_1882) | (n_3343 & n_1881));
 assign n_3364 = ((n_2833 & n_1885) | (n_3344 & n_1881));
 assign n_3365 = ((n_2833 & n_1888) | (n_3345 & n_1881));
 assign n_3366 = ((n_2833 & n_1889) | (n_3347 & n_1881));
 assign n_3367 = ((n_2833 & n_1896) | (n_3348 & n_1881));
 assign n_3368 = ((n_2833 & n_1897) | (n_3349 & n_1881));
 assign n_3369 = ((n_2833 & n_1886) | (n_3350 & n_1881));
 assign n_3370 = ((n_2833 & n_1890) | (n_3351 & n_1881));
 assign n_3371 = ((n_2833 & n_1898) | (n_3352 & n_1881));
 assign n_3372 = ((n_2833 & n_1901) | (n_3358 & n_1881));
 assign n_3373 = ((n_2833 & n_1891) | (n_3354 & n_1881));
 assign n_3374 = ((n_2833 & n_1883) | (n_3356 & n_1881));
 assign n_3375 = ((n_2833 & n_1884) | (n_3357 & n_1881));
 assign n_3376 = ((n_2833 & n_1899) | (n_3353 & n_1881));
 assign n_3377 = ((n_2833 & n_493) | (n_1881 & n_496));
 assign n_3378 = ((n_2833 & n_1887) | (n_3359 & n_1881));
 assign n_3379 = ((n_2833 & n_1892) | (n_3360 & n_1881));
 assign n_3380 = ((n_2833 & n_1893) | (n_3361 & n_1881));
 assign n_3381 = ((n_2833 & n_1894) | (n_3362 & n_1881));
 assign n_3382 = ((n_2863 & n_880) | (n_882 & n_1924));
 assign n_3383 = ((n_2863 & n_1928) | (n_888 & n_1924));
 assign n_3384 = ((n_2863 & n_1931) | (n_909 & n_1924));
 assign n_3385 = ((n_2863 & n_884) | (n_889 & n_1924));
 assign n_3386 = ((n_2863 & n_1932) | (n_911 & n_1924));
 assign n_3387 = ((n_2863 & n_1925) | (n_912 & n_1924));
 assign n_3388 = ((n_2863 & n_879) | (n_881 & n_1924));
 assign n_3389 = ((n_2863 & n_1929) | (n_878 & n_1924));
 assign n_3390 = ((n_2863 & n_3705) | (n_877 & n_1924));
 assign n_3391 = ((n_2863 & n_871) | (n_872 & n_1924));
 assign n_3392 = ((n_2863 & n_868) | (n_864 & n_1924));
 assign n_3393 = ((n_2863 & n_854) | (n_855 & n_1924));
 assign n_3394 = ((n_2863 & n_869) | (n_866 & n_1924));
 assign n_3395 = ((n_2863 & n_1926) | (n_865 & n_1924));
 assign n_3396 = ((n_2863 & n_1927) | (n_902 & n_1924));
 assign n_3397 = ((n_2863 & n_867) | (n_870 & n_1924));
 assign n_3398 = ((n_2863 & n_1934) | (n_900 & n_1924));
 assign n_3399 = ((n_2863 & n_1930) | (n_861 & n_1924));
 assign n_3400 = ((n_2863 & n_1935) | (n_860 & n_1924));
 assign n_3401 = ((n_2863 & n_672) | (n_1924 & n_710));
 assign n_3402 = ((n_2863 & n_896) | (n_901 & n_1924));
 assign n_3403 = ((n_2863 & n_883) | (n_856 & n_1924));
 assign n_3404 = ((n_2889 & n_1984) | (n_3382 & n_1969));
 assign n_3405 = ((n_2889 & n_1973) | (n_3383 & n_1969));
 assign n_3406 = ((n_2889 & n_1976) | (n_3384 & n_1969));
 assign n_3407 = ((n_2889 & n_1983) | (n_3385 & n_1969));
 assign n_3408 = ((n_2889 & n_1977) | (n_3386 & n_1969));
 assign n_3409 = ((n_2889 & n_1970) | (n_3387 & n_1969));
 assign n_3410 = ((n_2889 & n_1985) | (n_3388 & n_1969));
 assign n_3411 = ((n_2889 & n_1974) | (n_3389 & n_1969));
 assign n_3412 = ((n_2889 & n_1978) | (n_3390 & n_1969));
 assign n_3413 = ((n_2889 & n_1986) | (n_3391 & n_1969));
 assign n_3414 = ((n_2889 & n_1987) | (n_3392 & n_1969));
 assign n_3415 = ((n_2889 & n_1975) | (n_3399 & n_1969));
 assign n_3416 = ((n_2889 & n_1988) | (n_3394 & n_1969));
 assign n_3417 = ((n_2889 & n_1971) | (n_3395 & n_1969));
 assign n_3418 = ((n_2889 & n_1972) | (n_3396 & n_1969));
 assign n_3419 = ((n_2889 & n_1989) | (n_3397 & n_1969));
 assign n_3420 = ((n_2889 & n_1990) | (n_3393 & n_1969));
 assign n_3421 = ((n_2889 & n_1979) | (n_3398 & n_1969));
 assign n_3422 = ((n_2889 & n_1980) | (n_3400 & n_1969));
 assign n_3423 = ((n_2889 & n_1991) | (n_3401 & n_1969));
 assign n_3424 = ((n_2889 & n_1981) | (n_3402 & n_1969));
 assign n_3425 = ((n_2889 & n_569) | (n_1969 & n_574));
 assign n_3426 = ((n_2889 & n_1982) | (n_3403 & n_1969));
 assign n_3427 = ((n_300 & n_2032) | (n_3410 & n_2016));
 assign n_3428 = ((n_300 & n_2020) | (n_3405 & n_2016));
 assign n_3429 = ((n_300 & n_2023) | (n_3406 & n_2016));
 assign n_3430 = ((n_300 & n_2030) | (n_3407 & n_2016));
 assign n_3431 = ((n_300 & n_2024) | (n_3408 & n_2016));
 assign n_3432 = ((n_300 & n_2031) | (n_3404 & n_2016));
 assign n_3433 = ((n_300 & n_2021) | (n_3411 & n_2016));
 assign n_3434 = ((n_300 & n_2025) | (n_3412 & n_2016));
 assign n_3435 = ((n_300 & n_2033) | (n_3413 & n_2016));
 assign n_3436 = ((n_300 & n_2034) | (n_3414 & n_2016));
 assign n_3437 = ((n_300 & n_2026) | (n_3421 & n_2016));
 assign n_3438 = ((n_300 & n_2027) | (n_3422 & n_2016));
 assign n_3439 = ((n_300 & n_2018) | (n_3417 & n_2016));
 assign n_3440 = ((n_300 & n_2019) | (n_3418 & n_2016));
 assign n_3441 = ((n_300 & n_2036) | (n_3419 & n_2016));
 assign n_3442 = ((n_300 & n_2037) | (n_3420 & n_2016));
 assign n_3443 = ((n_300 & n_2022) | (n_3415 & n_2016));
 assign n_3444 = ((n_300 & n_2035) | (n_3416 & n_2016));
 assign n_3445 = ((n_300 & n_2038) | (n_3423 & n_2016));
 assign n_3446 = ((n_300 & n_2028) | (n_3424 & n_2016));
 assign n_3447 = ((n_300 & n_2039) | (n_3425 & n_2016));
 assign n_3448 = ((n_300 & n_2029) | (n_3426 & n_2016));
 assign n_3449 = ((n_2949 & n_2081) | (n_916 & n_2065));
 assign n_3450 = ((n_2949 & n_2069) | (n_923 & n_2065));
 assign n_3451 = ((n_2949 & n_2072) | (n_924 & n_2065));
 assign n_3452 = ((n_2949 & n_2079) | (n_936 & n_2065));
 assign n_3453 = ((n_2949 & n_2073) | (n_925 & n_2065));
 assign n_3454 = ((n_2949 & n_3709) | (n_2041 & n_2065));
 assign n_3455 = ((n_2949 & n_2070) | (n_932 & n_2065));
 assign n_3456 = ((n_2949 & n_2074) | (n_922 & n_2065));
 assign n_3457 = ((n_2949 & n_2082) | (n_915 & n_2065));
 assign n_3458 = ((n_2949 & n_2075) | (n_919 & n_2065));
 assign n_3459 = ((n_2949 & n_2084) | (n_927 & n_2065));
 assign n_3460 = ((n_2949 & n_2067) | (n_914 & n_2065));
 assign n_3461 = ((n_2949 & n_2068) | (n_930 & n_2065));
 assign n_3462 = ((n_2949 & n_2085) | (n_935 & n_2065));
 assign n_3463 = ((n_2949 & n_2086) | (n_928 & n_2065));
 assign n_3464 = ((n_2949 & n_2071) | (n_934 & n_2065));
 assign n_3465 = ((n_2949 & n_2076) | (n_929 & n_2065));
 assign n_3466 = ((n_2949 & n_2087) | (n_918 & n_2065));
 assign n_3467 = ((n_2949 & n_2077) | (n_920 & n_2065));
 assign n_3468 = ((n_2949 & n_2088) | (n_917 & n_2065));
 assign n_3469 = ((n_2949 & n_2078) | (n_937 & n_2065));
 assign n_3470 = ((n_2979 & n_2117) | (n_3454 & n_2116));
 assign n_3471 = ((n_2979 & n_2120) | (n_3450 & n_2116));
 assign n_3472 = ((n_2979 & n_2123) | (n_3451 & n_2116));
 assign n_3473 = ((n_2979 & n_2130) | (n_3452 & n_2116));
 assign n_3474 = ((n_2979 & n_2124) | (n_3453 & n_2116));
 assign n_3475 = ((n_2979 & n_2131) | (n_2105 & n_2116));
 assign n_3476 = ((n_2979 & n_2132) | (n_3449 & n_2116));
 assign n_3477 = ((n_2979 & n_2121) | (n_3455 & n_2116));
 assign n_3478 = ((n_2979 & n_2125) | (n_3456 & n_2116));
 assign n_3479 = ((n_2979 & n_2133) | (n_3457 & n_2116));
 assign n_3480 = ((n_2979 & n_2126) | (n_3458 & n_2116));
 assign n_3481 = ((n_2979 & n_2135) | (n_3459 & n_2116));
 assign n_3482 = ((n_2979 & n_2118) | (n_3460 & n_2116));
 assign n_3483 = ((n_2979 & n_2119) | (n_3461 & n_2116));
 assign n_3484 = ((n_2979 & n_2136) | (n_3462 & n_2116));
 assign n_3485 = ((n_2979 & n_2137) | (n_3463 & n_2116));
 assign n_3486 = ((n_2979 & n_2122) | (n_3464 & n_2116));
 assign n_3487 = ((n_2979 & n_2127) | (n_3465 & n_2116));
 assign n_3488 = ((n_2979 & n_2138) | (n_3466 & n_2116));
 assign n_3489 = ((n_2979 & n_2128) | (n_3467 & n_2116));
 assign n_3490 = ((n_2979 & n_2139) | (n_3468 & n_2116));
 assign n_3491 = ((n_2979 & n_2129) | (n_3469 & n_2116));
 assign n_3492 = ((n_3009 & n_2170) | (n_992 & n_2169));
 assign n_3493 = ((n_3009 & n_2173) | (n_971 & n_2169));
 assign n_3494 = ((n_3009 & n_2176) | (n_964 & n_2169));
 assign n_3495 = ((n_3009 & n_2183) | (n_1006 & n_2169));
 assign n_3496 = ((n_3009 & n_2177) | (n_981 & n_2169));
 assign n_3497 = ((n_3009 & n_2184) | (n_1008 & n_2169));
 assign n_3498 = ((n_3009 & n_2185) | (n_994 & n_2169));
 assign n_3499 = ((n_3009 & n_2174) | (n_945 & n_2169));
 assign n_3500 = ((n_3009 & n_2178) | (n_1009 & n_2169));
 assign n_3501 = ((n_3009 & n_2186) | (n_984 & n_2169));
 assign n_3502 = ((n_3009 & n_1001) | (n_955 & n_2169));
 assign n_3503 = ((n_3009 & n_2179) | (n_1012 & n_2169));
 assign n_3504 = ((n_3009 & n_2171) | (n_975 & n_2169));
 assign n_3505 = ((n_3009 & n_2172) | (n_963 & n_2169));
 assign n_3506 = ((n_3009 & n_969) | (n_939 & n_2169));
 assign n_3507 = ((n_3009 & n_2175) | (n_954 & n_2169));
 assign n_3508 = ((n_3009 & n_2180) | (n_1014 & n_2169));
 assign n_3509 = ((n_3009 & n_968) | (n_972 & n_2169));
 assign n_3510 = ((n_3009 & n_2181) | (n_988 & n_2169));
 assign n_3511 = ((n_3009 & n_956) | (n_941 & n_2169));
 assign n_3512 = ((n_3009 & n_2182) | (n_949 & n_2169));
 assign n_3513 = ((n_3009 & n_958) | (n_948 & n_2169));
 assign n_3514 = ((n_3009 & n_1000) | (n_985 & n_2169));
 assign n_3515 = ((n_3034 & n_2234) | (n_3503 & n_2224));
 assign n_3516 = ((n_3034 & n_2238) | (n_3495 & n_2224));
 assign n_3517 = ((n_3034 & n_379) | (n_2224 & n_366));
 assign n_3518 = ((n_3034 & n_2239) | (n_3497 & n_2224));
 assign n_3519 = ((n_3034 & n_2240) | (n_3498 & n_2224));
 assign n_3520 = ((n_3034 & n_2229) | (n_3499 & n_2224));
 assign n_3521 = ((n_3034 & n_2233) | (n_3500 & n_2224));
 assign n_3522 = ((n_3034 & n_2241) | (n_3501 & n_2224));
 assign n_3523 = ((n_3034 & n_2242) | (n_3502 & n_2224));
 assign n_3524 = ((n_3034 & n_2225) | (n_3492 & n_2224));
 assign n_3525 = ((n_3034 & n_2250) | (n_3065 & n_2224));
 assign n_3526 = ((n_3034 & n_2244) | (n_3066 & n_2224));
 assign n_3527 = ((n_3034 & n_2245) | (n_3506 & n_2224));
 assign n_3528 = ((n_3034 & n_2235) | (n_3508 & n_2224));
 assign n_3529 = ((n_3034 & n_2246) | (n_3509 & n_2224));
 assign n_3530 = ((n_3034 & n_2236) | (n_3510 & n_2224));
 assign n_3531 = ((n_3034 & n_2247) | (n_3511 & n_2224));
 assign n_3532 = ((n_3034 & n_2248) | (n_3067 & n_2224));
 assign n_3533 = ((n_3034 & n_2237) | (n_3512 & n_2224));
 assign n_3534 = ((n_3034 & n_2249) | (n_3513 & n_2224));
 assign n_3535 = ((n_3034 & n_2243) | (n_3514 & n_2224));
 assign n_3536 = ~(sub_181_2_n_0 & (~{in2[30]} | {in1[0]}));
 assign n_3537 = ~({in1[24]} | ({in1[25]} | (~n_3105 | ~n_3102)));
 assign n_3538 = (n_3183 & (sub_219_2_n_37 | sub_219_2_n_9));
 assign n_3540 = (~sub_276_2_n_6 & (n_3234 | sub_276_2_n_13));
 assign n_3541 = (~sub_276_2_n_0 & (sub_276_2_n_7 | sub_276_2_n_18));
 assign n_3542 = (sub_295_2_n_1 & (sub_295_2_n_22 | sub_295_2_n_10));
 assign n_3543 = ~(sub_314_2_n_3 & (sub_314_2_n_37 & (sub_314_2_n_30 & ~n_401)));
 assign n_3544 = ((n_741 & n_740) | (n_748 & n_736));
 assign n_3545 = (sub_352_2_n_29 & (sub_352_2_n_63 | sub_352_2_n_27));
 assign n_3546 = (sub_352_2_n_32 & (n_3176 | sub_352_2_n_20));
 assign n_3547 = ~(sub_371_2_n_9 | (~sub_371_2_n_19 | ~n_3251));
 assign n_3548 = (~sub_371_2_n_9 & (n_3251 | sub_371_2_n_19));
 assign n_3549 = ~(sub_390_2_n_95 & (sub_390_2_n_69 & (~sub_390_2_n_76 & ~n_354)));
 assign n_3550 = (sub_390_2_n_1 | (sub_390_2_n_96 & sub_390_2_n_53));
 assign n_3551 = ~((~sub_390_2_n_47 | ~sub_390_2_n_50) & (sub_390_2_n_74 | sub_390_2_n_70));
 assign n_3552 = (~n_3204 | (sub_390_2_n_71 & sub_390_2_n_96));
 assign n_3553 = ~(sub_409_2_n_23 & (~n_3175 | sub_409_2_n_51));
 assign n_3554 = (~sub_409_2_n_71 | (sub_409_2_n_68 & n_3175));
 assign n_3555 = ~(n_3174 & (~sub_409_2_n_101 | sub_409_2_n_52));
 assign n_3556 = ~(sub_428_2_n_57 & (~sub_428_2_n_103 | sub_428_2_n_56));
 assign n_3557 = (sub_428_2_n_4 & (sub_428_2_n_85 | sub_428_2_n_30));
 assign n_3558 = ~((~sub_428_2_n_58 | ~sub_428_2_n_47) & (sub_428_2_n_78 | sub_428_2_n_74));
 assign n_3559 = (~sub_428_2_n_34 & (n_3276 | sub_428_2_n_41));
 assign n_3560 = (~sub_428_2_n_80 | (n_3559 & sub_428_2_n_103));
 assign n_3561 = ~(sub_428_2_n_78 & (~sub_428_2_n_95 | sub_428_2_n_14));
 assign n_3562 = (~sub_428_2_n_8 | (sub_428_2_n_95 & sub_428_2_n_29));
 assign n_3563 = ~((~sub_447_2_n_88 & ~sub_447_2_n_76) | (sub_447_2_n_3 & sub_447_2_n_60));
 assign n_3564 = (sub_447_2_n_5 & (sub_447_2_n_26 | sub_447_2_n_28));
 assign n_3565 = ~(n_793 & (~n_3171 | n_792));
 assign n_3566 = ~(n_822 & (~sub_466_2_n_107 | n_824));
 assign n_3567 = (~n_817 | (n_813 & n_3171));
 assign n_3568 = (~n_831 | (n_830 & sub_466_2_n_122));
 assign n_3569 = (~sub_485_2_n_0 | (sub_485_2_n_110 & sub_485_2_n_48));
 assign n_3570 = ~(sub_485_2_n_8 & (~sub_485_2_n_37 | n_3210));
 assign n_3571 = ~(sub_485_2_n_95 | (~sub_485_2_n_85 | ~n_3144));
 assign n_3572 = ~((~sub_485_2_n_0 & ~sub_485_2_n_55) | (sub_485_2_n_82 & sub_485_2_n_79));
 assign n_3573 = (sub_485_2_n_2 & (sub_485_2_n_49 | sub_485_2_n_51));
 assign n_3574 = (~sub_504_2_n_88 | (sub_504_2_n_71 & sub_504_2_n_121));
 assign n_3575 = ~(n_3586 & (~sub_504_2_n_129 | sub_504_2_n_67));
 assign n_3576 = (~sub_504_2_n_55 | (sub_504_2_n_129 & sub_504_2_n_9));
 assign n_3577 = (~n_3587 | (sub_504_2_n_128 & sub_504_2_n_83));
 assign n_3578 = (~sub_504_2_n_52 | (sub_504_2_n_128 & sub_504_2_n_37));
 assign n_3579 = (~sub_504_2_n_38 | (n_3574 & sub_504_2_n_31));
 assign n_3580 = ~(sub_504_2_n_34 & (~sub_504_2_n_121 | sub_504_2_n_32));
 assign n_3581 = (~sub_504_2_n_44 | (n_3582 & sub_504_2_n_45));
 assign n_3582 = ~(sub_504_2_n_86 & (~sub_504_2_n_109 | sub_504_2_n_84));
 assign n_3583 = (~sub_504_2_n_7 | (sub_504_2_n_109 & sub_504_2_n_5));
 assign n_3584 = (sub_504_2_n_1 | (sub_504_2_n_101 & sub_504_2_n_51));
 assign n_3585 = ((n_3586 | sub_504_2_n_81) & (sub_504_2_n_47 | n_453));
 assign n_3586 = (~sub_504_2_n_8 & (sub_504_2_n_55 | sub_504_2_n_56));
 assign n_3587 = (sub_504_2_n_0 & (sub_504_2_n_52 | sub_504_2_n_53));
 assign n_3588 = (~sub_523_2_n_40 | (sub_523_2_n_27 & sub_523_2_n_57));
 assign n_3589 = (~sub_523_2_n_49 | (sub_523_2_n_131 & sub_523_2_n_44));
 assign n_3591 = (~sub_523_2_n_61 & (n_3592 | sub_523_2_n_53));
 assign n_3592 = (sub_523_2_n_101 & (sub_523_2_n_123 | sub_523_2_n_95));
 assign n_3593 = (~sub_523_2_n_46 | (n_3596 & sub_523_2_n_37));
 assign n_3594 = (sub_523_2_n_54 | (n_840 & sub_523_2_n_41));
 assign n_3595 = ~((~sub_523_2_n_0 & ~sub_523_2_n_62) | (sub_523_2_n_91 & sub_523_2_n_88));
 assign n_3596 = ~(sub_523_2_n_89 & (~n_3701 | sub_523_2_n_22));
 assign n_3597 = (~sub_542_2_n_47 | (sub_542_2_n_135 & sub_542_2_n_0));
 assign n_3598 = (~sub_542_2_n_43 | (n_3602 & sub_542_2_n_13));
 assign n_3599 = ~(n_3607 & (~n_3602 | sub_542_2_n_94));
 assign n_3600 = ~(sub_542_2_n_110 | (sub_542_2_n_102 | n_3692));
 assign n_3601 = (~sub_542_2_n_53 | (sub_542_2_n_137 & sub_542_2_n_4));
 assign n_3602 = (sub_542_2_n_24 | (sub_542_2_n_103 & sub_542_2_n_129));
 assign n_3603 = (~sub_542_2_n_42 | (sub_542_2_n_129 & sub_542_2_n_2));
 assign n_3604 = ~(sub_542_2_n_103 & (sub_542_2_n_104 & sub_542_2_n_129));
 assign n_3605 = (~sub_542_2_n_3 | (n_3703 & sub_542_2_n_58));
 assign n_3606 = (sub_542_2_n_6 | (sub_542_2_n_113 & sub_542_2_n_62));
 assign n_3607 = (sub_542_2_n_67 & (sub_542_2_n_43 | sub_542_2_n_55));
 assign n_3608 = (sub_542_2_n_11 | (n_3599 & sub_542_2_n_64));
 assign n_3609 = (~n_862 | (n_3611 & n_863));
 assign n_3610 = (~n_887 | (n_3612 & n_885));
 assign n_3611 = (~n_891 | (n_906 & n_893));
 assign n_3612 = ~(n_874 & (~n_906 | n_875));
 assign n_3613 = (~n_857 | (n_906 & n_859));
 assign n_3614 = ~(sub_561_2_n_145 & (sub_561_2_n_72 & (n_3619 & ~sub_561_2_n_119)));
 assign n_3615 = (sub_561_2_n_117 & (sub_561_2_n_138 | sub_561_2_n_109));
 assign n_3616 = (~sub_561_2_n_2 | (n_3707 & sub_561_2_n_6));
 assign n_3617 = (sub_561_2_n_11 | (sub_561_2_n_121 & sub_561_2_n_62));
 assign n_3618 = (n_3620 & (n_3621 | sub_561_2_n_100));
 assign n_3619 = ~((~sub_561_2_n_0 & ~sub_561_2_n_40) | (sub_561_2_n_105 & sub_561_2_n_98));
 assign n_3620 = (sub_561_2_n_70 & (sub_561_2_n_63 | sub_561_2_n_50));
 assign n_3621 = ~(sub_561_2_n_73 | (~sub_561_2_n_39 & sub_561_2_n_41));
 assign n_3622 = (~sub_580_2_n_104 | (sub_580_2_n_98 & sub_580_2_n_153));
 assign n_3623 = ~(sub_580_2_n_2 & (~sub_580_2_n_153 | sub_580_2_n_66));
 assign n_3624 = ~(sub_580_2_n_49 & (~n_3626 | sub_580_2_n_77));
 assign n_3625 = (~sub_580_2_n_11 | (n_3628 & sub_580_2_n_68));
 assign n_3626 = (~sub_580_2_n_24 | (sub_580_2_n_99 & sub_580_2_n_140));
 assign n_3627 = ~(sub_580_2_n_56 & (~sub_580_2_n_140 | sub_580_2_n_47));
 assign n_3628 = (sub_580_2_n_102 | (sub_580_2_n_94 & sub_580_2_n_139));
 assign n_3629 = (~sub_580_2_n_9 | (sub_580_2_n_139 & sub_580_2_n_75));
 assign n_3630 = (~sub_580_2_n_15 | (sub_580_2_n_131 & sub_580_2_n_55));
 assign n_3631 = (sub_580_2_n_44 | (sub_580_2_n_117 & sub_580_2_n_69));
 assign n_3632 = ~((~sub_580_2_n_11 & ~sub_580_2_n_73) | (sub_580_2_n_102 & sub_580_2_n_97));
 assign n_3633 = (sub_599_2_n_129 & (sub_599_2_n_145 | sub_599_2_n_122));
 assign n_3634 = ~(sub_599_2_n_14 & (~sub_599_2_n_141 | sub_599_2_n_69));
 assign n_3635 = ~((~sub_599_2_n_14 & ~sub_599_2_n_62) | (sub_599_2_n_111 & sub_599_2_n_95));
 assign n_3636 = ~((~sub_599_2_n_73 & ~sub_599_2_n_77) | (sub_599_2_n_117 & sub_599_2_n_107));
 assign n_3637 = (~sub_618_2_n_7 | (n_3638 & sub_618_2_n_0));
 assign n_3638 = ~(sub_618_2_n_25 & (~sub_618_2_n_174 | sub_618_2_n_110));
 assign n_3639 = (~sub_618_2_n_69 | (sub_618_2_n_174 & sub_618_2_n_2));
 assign n_3640 = (~sub_618_2_n_81 | (n_3652 & sub_618_2_n_50));
 assign n_3641 = (~sub_618_2_n_82 | (n_3654 & sub_618_2_n_64));
 assign n_3642 = (~sub_618_2_n_6 | (sub_618_2_n_161 & sub_618_2_n_76));
 assign n_3643 = (~sub_618_2_n_1 | (n_3645 & sub_618_2_n_56));
 assign n_3644 = ~(sub_618_2_n_11 & (~n_3647 | sub_618_2_n_78));
 assign n_3645 = (sub_618_2_n_116 | (sub_618_2_n_107 & sub_618_2_n_152));
 assign n_3646 = (~sub_618_2_n_77 | (sub_618_2_n_152 & sub_618_2_n_54));
 assign n_3647 = ~(sub_618_2_n_130 & (~sub_618_2_n_152 | sub_618_2_n_120));
 assign n_3648 = (~sub_618_2_n_14 | (n_3653 & sub_618_2_n_60));
 assign n_3649 = (~sub_618_2_n_12 | (sub_618_2_n_142 & sub_618_2_n_8));
 assign n_3650 = ~((~sub_618_2_n_82 & ~sub_618_2_n_70) | (sub_618_2_n_117 & sub_618_2_n_108));
 assign n_3651 = ~(sub_618_2_n_68 | (n_3154 | (~sub_618_2_n_42 | ~n_3153)));
 assign n_3652 = (~sub_618_2_n_121 | (sub_618_2_n_113 & sub_618_2_n_161));
 assign n_3653 = ~(sub_618_2_n_118 & (~sub_618_2_n_142 | sub_618_2_n_109));
 assign n_3654 = (sub_618_2_n_117 | (sub_618_2_n_111 & n_3647));
 assign n_3655 = ~(n_3153 & (sub_618_2_n_42 & (~sub_618_2_n_66 & ~n_3154)));
 assign n_3656 = (~sub_637_2_n_64 | (sub_637_2_n_189 & sub_637_2_n_55));
 assign n_3657 = (~sub_637_2_n_68 | (sub_637_2_n_175 & sub_637_2_n_41));
 assign n_3658 = (~sub_637_2_n_72 | (sub_637_2_n_173 & sub_637_2_n_9));
 assign n_3659 = (~sub_637_2_n_63 | (sub_637_2_n_163 & sub_637_2_n_48));
 assign n_3660 = (~sub_637_2_n_74 | (sub_637_2_n_150 & sub_637_2_n_52));
 assign n_3661 = (sub_637_2_n_116 & (sub_637_2_n_119 | sub_637_2_n_16));
 assign n_3662 = ~((~sub_637_2_n_5 & ~sub_637_2_n_42) | (sub_637_2_n_123 & sub_637_2_n_96));
 assign n_3663 = ~((~sub_637_2_n_64 & ~sub_637_2_n_73) | (sub_637_2_n_121 & sub_637_2_n_114));
 assign n_3664 = ~(sub_637_2_n_40 | (sub_637_2_n_45 | (~sub_637_2_n_94 | ~n_3153)));
 assign n_3665 = (~sub_637_2_n_4 & (sub_637_2_n_56 | sub_637_2_n_43));
 assign n_3666 = ~(sub_637_2_n_135 | (~sub_637_2_n_158 & sub_637_2_n_125));
 assign n_3667 = ~(n_967 & (~n_1002 | n_976));
 assign n_3668 = (~n_940 | (n_3670 & n_942));
 assign n_3669 = ~(n_1015 & (~n_3667 | n_966));
 assign n_3670 = (~n_952 | (n_951 & n_3673));
 assign n_3671 = ~(n_944 & (~n_3673 | n_943));
 assign n_3672 = ~(n_962 & (~n_3674 | n_1005));
 assign n_3673 = (~n_1004 | (n_1002 & n_978));
 assign n_3674 = ~(n_986 & (~n_1002 | n_1010));
 assign n_3675 = (~n_1013 | (n_1002 & n_980));
 assign n_3676 = (~n_983 | (n_977 & n_982));
 assign n_3677 = (~sub_656_2_n_128 | (sub_656_2_n_99 & sub_656_2_n_157));
 assign n_3678 = (~sub_656_2_n_78 | (n_3748 & sub_656_2_n_39));
 assign n_3679 = (~sub_675_2_n_68 | (n_3680 & sub_675_2_n_39));
 assign n_3680 = (~n_3684 | (sub_675_2_n_116 & sub_675_2_n_169));
 assign n_3681 = ~(sub_675_2_n_139 & (~n_3177 | sub_675_2_n_129));
 assign n_3682 = ~((~sub_675_2_n_1 & ~sub_675_2_n_47) | (sub_675_2_n_125 & sub_675_2_n_96));
 assign n_3683 = (sub_675_2_n_12 & (sub_675_2_n_68 | sub_675_2_n_46));
 assign n_3684 = (~sub_675_2_n_6 & (sub_675_2_n_40 | sub_675_2_n_33));
 assign n_3685 = (~sub_675_2_n_72 & (sub_675_2_n_60 | sub_675_2_n_59));
 assign n_3686 = (~sub_694_2_n_143 & (sub_694_2_n_169 | sub_694_2_n_124));
 assign n_3687 = ((sub_694_2_n_136 | sub_694_2_n_124) & (sub_694_2_n_129 | sub_694_2_n_119));
 assign n_3688 = ~((sub_694_2_n_51 | sub_694_2_n_48) & (sub_694_2_n_114 | sub_694_2_n_106));
 assign n_3689 = ~(n_3113 & (~{in1[4]} & ~{in1[5]}));
 assign n_3690 = ~({in1[18]} | ({in1[19]} | (~n_3717 | ~n_3716)));
 assign n_3692 = ~(sub_542_2_n_135 & (~sub_542_2_n_93 & ~sub_542_2_n_19));
 assign n_3693 = ~((n_300 & n_512) | (n_2016 & n_514));
 assign n_3695 = (sub_447_2_n_64 & ~(sub_447_2_n_100 & n_3694));
 assign n_3694 = ~(~n_3288 & n_423);
 assign n_3697 = (sub_466_2_n_80 ^ n_3696);
 assign n_3696 = ~(n_797 | (~n_784 & n_3568));
 assign n_3699 = ~(sub_523_2_n_112 | (n_3749 & sub_523_2_n_131));
 assign n_3701 = ~(~sub_523_2_n_6 & (sub_523_2_n_65 | n_3700));
 assign n_3700 = ~(sub_523_2_n_54 | (sub_523_2_n_41 & n_840));
 assign n_3703 = ~(~sub_542_2_n_12 & (sub_542_2_n_69 | n_3702));
 assign n_3702 = ~(sub_542_2_n_6 | (sub_542_2_n_62 & sub_542_2_n_113));
 assign n_3705 = ~(n_876 ^ n_3704);
 assign n_3704 = ~(n_899 & (~n_895 | n_894));
 assign n_3707 = ~(~sub_561_2_n_1 & (sub_561_2_n_68 | n_3706));
 assign n_3706 = ~(sub_561_2_n_11 | (sub_561_2_n_121 & sub_561_2_n_62));
 assign n_3709 = ~(sub_618_2_n_24 ^ n_3708);
 assign n_3708 = ~(sub_618_2_n_136 | (~sub_618_2_n_126 & sub_618_2_n_161));
 assign n_3711 = ~(n_3710 & (~sub_656_2_n_26 | sub_656_2_n_130));
 assign n_3710 = ~(~sub_656_2_n_165 | (sub_656_2_n_12 | sub_656_2_n_23));
 assign n_3713 = ~(sub_447_2_n_25 & (~n_3207 | n_3712));
 assign n_3712 = (sub_447_2_n_64 & (sub_447_2_n_97 | sub_447_2_n_46));
 assign n_3715 = ~(n_3083 & (n_3080 & n_3714));
 assign n_3714 = ~({in1[12]} | ({in1[13]} | ~n_3690));
 assign n_3716 = ~({in1[16]} | {in1[17]});
 assign n_3717 = ~({in1[14]} | {in1[15]});
 assign n_3718 = ~({in1[30]} | {in1[31]});
 assign n_3719 = ~(n_3095 & (n_3092 & n_3718));
 assign n_3720 = ~(n_3159 | n_3719);
 assign n_3721 = ((n_1507 & n_2567) | (n_3227 & n_1504));
 assign n_3722 = ((n_1506 & n_2567) | (n_3239 & n_1504));
 assign n_3723 = ((n_1509 & n_2567) | (n_3240 & n_1504));
 assign n_3724 = ((n_1510 & n_2567) | (n_1502 & n_1504));
 assign n_3725 = ((n_1566 & n_2607) | (n_3246 & n_1561));
 assign n_3726 = ((n_1570 & n_2607) | (n_3248 & n_1561));
 assign n_3727 = ((n_1571 & n_2607) | (n_3038 & n_1561));
 assign n_3728 = ((n_2719 & n_1743) | (n_812 & n_1729));
 assign n_3729 = ((n_2719 & n_1730) | (n_806 & n_1729));
 assign n_3730 = ((n_2719 & n_1742) | (n_809 & n_1729));
 assign n_3731 = ((n_2719 & n_3697) | (n_800 & n_1729));
 assign n_3732 = ((n_2747 & n_1771) | (n_3309 & n_2748));
 assign n_3733 = ((n_1772 & n_2747) | (n_3307 & n_2748));
 assign n_3734 = ((n_2747 & n_1779) | (n_3055 & n_1764));
 assign n_3735 = ((n_2781 & n_1810) | (n_1791 & n_1801));
 assign n_3736 = ((n_2781 & n_1805) | (n_3321 & n_1801));
 assign n_3737 = ((n_2781 & n_1808) | (n_3732 & n_1801));
 assign n_3738 = ((n_2781 & n_1815) | (n_3322 & n_1801));
 assign n_3739 = ((n_2781 & n_1816) | (n_3734 & n_1801));
 assign n_3740 = ((n_2781 & n_1818) | (n_1799 & n_1801));
 assign n_3741 = ((n_2781 & n_1819) | (n_3058 & n_1801));
 assign n_3742 = ((n_2781 & n_1811) | (n_3326 & n_1801));
 assign n_3743 = ((n_2781 & n_1812) | (n_3329 & n_1801));
 assign n_3744 = ((n_2781 & n_1814) | (n_3325 & n_1801));
 assign n_3745 = (~sub_409_2_n_3 | (n_3554 & sub_409_2_n_49));
 assign n_3746 = (sub_428_2_n_9 & (n_3182 | sub_428_2_n_48));
 assign n_3747 = (~sub_656_2_n_42 | (sub_656_2_n_157 & sub_656_2_n_51));
 assign n_3748 = ~(sub_656_2_n_125 & (~sub_656_2_n_148 | sub_656_2_n_17));
 assign n_3749 = (sub_523_2_n_75 & (sub_523_2_n_74 & (sub_523_2_n_102 & sub_523_2_n_87)));
endmodule


