`timescale 1ps / 1ps
module fft2_Mul_32Sx21S_50S_4(
          in2,
          in1,
          out1,
          clk,
          clr
);
   input [31:0] in2;
   input [20:0] in1;
   output [49:0] out1;
   input clk;
   input clr;
wire mul_22_25_n_0, mul_22_25_n_1, mul_22_25_n_2, mul_22_25_n_3, mul_22_25_n_4,
     mul_22_25_n_5, mul_22_25_n_6, mul_22_25_n_7, mul_22_25_n_8, mul_22_25_n_9,
     mul_22_25_n_11, mul_22_25_n_12, mul_22_25_n_13, mul_22_25_n_14,
     mul_22_25_n_15, mul_22_25_n_16, mul_22_25_n_19, mul_22_25_n_20,
     mul_22_25_n_21, mul_22_25_n_22, mul_22_25_n_23, mul_22_25_n_24,
     mul_22_25_n_25, mul_22_25_n_26, mul_22_25_n_27, mul_22_25_n_28,
     mul_22_25_n_29, mul_22_25_n_30, mul_22_25_n_31, mul_22_25_n_32,
     mul_22_25_n_33, mul_22_25_n_34, mul_22_25_n_35, mul_22_25_n_36,
     mul_22_25_n_37, mul_22_25_n_38, mul_22_25_n_39, mul_22_25_n_40,
     mul_22_25_n_41, mul_22_25_n_42, mul_22_25_n_43, mul_22_25_n_44,
     mul_22_25_n_45, mul_22_25_n_46, mul_22_25_n_47, mul_22_25_n_48,
     mul_22_25_n_49, mul_22_25_n_50, mul_22_25_n_51, mul_22_25_n_52,
     mul_22_25_n_53, mul_22_25_n_54, mul_22_25_n_55, mul_22_25_n_56,
     mul_22_25_n_57, mul_22_25_n_58, mul_22_25_n_59, mul_22_25_n_60,
     mul_22_25_n_61, mul_22_25_n_62, mul_22_25_n_63, mul_22_25_n_64,
     mul_22_25_n_65, mul_22_25_n_66, mul_22_25_n_67, mul_22_25_n_68,
     mul_22_25_n_69, mul_22_25_n_70, mul_22_25_n_71, mul_22_25_n_72,
     mul_22_25_n_73, mul_22_25_n_74, mul_22_25_n_75, mul_22_25_n_76,
     mul_22_25_n_77, mul_22_25_n_78, mul_22_25_n_79, mul_22_25_n_80,
     mul_22_25_n_81, mul_22_25_n_82, mul_22_25_n_83, mul_22_25_n_84,
     mul_22_25_n_85, mul_22_25_n_86, mul_22_25_n_87, mul_22_25_n_88,
     mul_22_25_n_89, mul_22_25_n_90, mul_22_25_n_91, mul_22_25_n_92,
     mul_22_25_n_94, mul_22_25_n_95, mul_22_25_n_96, mul_22_25_n_97,
     mul_22_25_n_98, mul_22_25_n_100, mul_22_25_n_101, mul_22_25_n_102,
     mul_22_25_n_103, mul_22_25_n_104, mul_22_25_n_105, mul_22_25_n_106,
     mul_22_25_n_107, mul_22_25_n_108, mul_22_25_n_109, mul_22_25_n_110,
     mul_22_25_n_111, mul_22_25_n_112, mul_22_25_n_113, mul_22_25_n_114,
     mul_22_25_n_115, mul_22_25_n_116, mul_22_25_n_117, mul_22_25_n_118,
     mul_22_25_n_119, mul_22_25_n_120, mul_22_25_n_121, mul_22_25_n_122,
     mul_22_25_n_123, mul_22_25_n_124, mul_22_25_n_125, mul_22_25_n_126,
     mul_22_25_n_127, mul_22_25_n_128, mul_22_25_n_129, mul_22_25_n_130,
     mul_22_25_n_131, mul_22_25_n_132, mul_22_25_n_133, mul_22_25_n_134,
     mul_22_25_n_135, mul_22_25_n_136, mul_22_25_n_137, mul_22_25_n_138,
     mul_22_25_n_139, mul_22_25_n_140, mul_22_25_n_141, mul_22_25_n_142,
     mul_22_25_n_143, mul_22_25_n_144, mul_22_25_n_145, mul_22_25_n_146,
     mul_22_25_n_147, mul_22_25_n_148, mul_22_25_n_149, mul_22_25_n_150,
     mul_22_25_n_151, mul_22_25_n_152, mul_22_25_n_153, mul_22_25_n_154,
     mul_22_25_n_155, mul_22_25_n_156, mul_22_25_n_157, mul_22_25_n_158,
     mul_22_25_n_159, mul_22_25_n_160, mul_22_25_n_161, mul_22_25_n_162,
     mul_22_25_n_163, mul_22_25_n_164, mul_22_25_n_165, mul_22_25_n_166,
     mul_22_25_n_167, mul_22_25_n_168, mul_22_25_n_169, mul_22_25_n_170,
     mul_22_25_n_171, mul_22_25_n_172, mul_22_25_n_173, mul_22_25_n_174,
     mul_22_25_n_175, mul_22_25_n_176, mul_22_25_n_177, mul_22_25_n_178,
     mul_22_25_n_179, mul_22_25_n_180, mul_22_25_n_181, mul_22_25_n_182,
     mul_22_25_n_183, mul_22_25_n_184, mul_22_25_n_185, mul_22_25_n_186,
     mul_22_25_n_187, mul_22_25_n_188, mul_22_25_n_189, mul_22_25_n_190,
     mul_22_25_n_191, mul_22_25_n_192, mul_22_25_n_193, mul_22_25_n_194,
     mul_22_25_n_195, mul_22_25_n_196, mul_22_25_n_197, mul_22_25_n_198,
     mul_22_25_n_199, mul_22_25_n_200, mul_22_25_n_201, mul_22_25_n_202,
     mul_22_25_n_203, mul_22_25_n_204, mul_22_25_n_205, mul_22_25_n_206,
     mul_22_25_n_207, mul_22_25_n_208, mul_22_25_n_209, mul_22_25_n_210,
     mul_22_25_n_211, mul_22_25_n_212, mul_22_25_n_213, mul_22_25_n_214,
     mul_22_25_n_215, mul_22_25_n_216, mul_22_25_n_217, mul_22_25_n_218,
     mul_22_25_n_219, mul_22_25_n_220, mul_22_25_n_221, mul_22_25_n_222,
     mul_22_25_n_223, mul_22_25_n_224, mul_22_25_n_225, mul_22_25_n_226,
     mul_22_25_n_227, mul_22_25_n_228, mul_22_25_n_229, mul_22_25_n_230,
     mul_22_25_n_231, mul_22_25_n_232, mul_22_25_n_233, mul_22_25_n_234,
     mul_22_25_n_235, mul_22_25_n_236, mul_22_25_n_237, mul_22_25_n_238,
     mul_22_25_n_239, mul_22_25_n_240, mul_22_25_n_241, mul_22_25_n_242,
     mul_22_25_n_243, mul_22_25_n_244, mul_22_25_n_245, mul_22_25_n_246,
     mul_22_25_n_247, mul_22_25_n_248, mul_22_25_n_249, mul_22_25_n_250,
     mul_22_25_n_251, mul_22_25_n_252, mul_22_25_n_253, mul_22_25_n_254,
     mul_22_25_n_255, mul_22_25_n_256, mul_22_25_n_257, mul_22_25_n_258,
     mul_22_25_n_259, mul_22_25_n_260, mul_22_25_n_261, mul_22_25_n_262,
     mul_22_25_n_263, mul_22_25_n_264, mul_22_25_n_265, mul_22_25_n_266,
     mul_22_25_n_267, mul_22_25_n_268, mul_22_25_n_269, mul_22_25_n_270,
     mul_22_25_n_271, mul_22_25_n_272, mul_22_25_n_273, mul_22_25_n_274,
     mul_22_25_n_275, mul_22_25_n_276, mul_22_25_n_277, mul_22_25_n_278,
     mul_22_25_n_279, mul_22_25_n_280, mul_22_25_n_281, mul_22_25_n_282,
     mul_22_25_n_283, mul_22_25_n_284, mul_22_25_n_285, mul_22_25_n_286,
     mul_22_25_n_287, mul_22_25_n_288, mul_22_25_n_289, mul_22_25_n_290,
     mul_22_25_n_291, mul_22_25_n_292, mul_22_25_n_293, mul_22_25_n_294,
     mul_22_25_n_295, mul_22_25_n_296, mul_22_25_n_297, mul_22_25_n_298,
     mul_22_25_n_299, mul_22_25_n_300, mul_22_25_n_301, mul_22_25_n_302,
     mul_22_25_n_303, mul_22_25_n_304, mul_22_25_n_305, mul_22_25_n_306,
     mul_22_25_n_307, mul_22_25_n_308, mul_22_25_n_309, mul_22_25_n_310,
     mul_22_25_n_311, mul_22_25_n_312, mul_22_25_n_313, mul_22_25_n_314,
     mul_22_25_n_315, mul_22_25_n_316, mul_22_25_n_317, mul_22_25_n_318,
     mul_22_25_n_319, mul_22_25_n_320, mul_22_25_n_321, mul_22_25_n_322,
     mul_22_25_n_323, mul_22_25_n_324, mul_22_25_n_325, mul_22_25_n_326,
     mul_22_25_n_327, mul_22_25_n_328, mul_22_25_n_329, mul_22_25_n_330,
     mul_22_25_n_331, mul_22_25_n_332, mul_22_25_n_333, mul_22_25_n_334,
     mul_22_25_n_335, mul_22_25_n_336, mul_22_25_n_337, mul_22_25_n_338,
     mul_22_25_n_339, mul_22_25_n_340, mul_22_25_n_341, mul_22_25_n_342,
     mul_22_25_n_343, mul_22_25_n_344, mul_22_25_n_345, mul_22_25_n_346,
     mul_22_25_n_347, mul_22_25_n_348, mul_22_25_n_349, mul_22_25_n_350,
     mul_22_25_n_351, mul_22_25_n_352, mul_22_25_n_353, mul_22_25_n_354,
     mul_22_25_n_355, mul_22_25_n_356, mul_22_25_n_357, mul_22_25_n_358,
     mul_22_25_n_359, mul_22_25_n_360, mul_22_25_n_361, mul_22_25_n_362,
     mul_22_25_n_363, mul_22_25_n_364, mul_22_25_n_365, mul_22_25_n_366,
     mul_22_25_n_367, mul_22_25_n_368, mul_22_25_n_369, mul_22_25_n_370,
     mul_22_25_n_371, mul_22_25_n_372, mul_22_25_n_373, mul_22_25_n_374,
     mul_22_25_n_375, mul_22_25_n_376, mul_22_25_n_377, mul_22_25_n_378,
     mul_22_25_n_379, mul_22_25_n_380, mul_22_25_n_381, mul_22_25_n_382,
     mul_22_25_n_383, mul_22_25_n_384, mul_22_25_n_385, mul_22_25_n_386,
     mul_22_25_n_387, mul_22_25_n_388, mul_22_25_n_389, mul_22_25_n_390,
     mul_22_25_n_391, mul_22_25_n_392, mul_22_25_n_393, mul_22_25_n_394,
     mul_22_25_n_395, mul_22_25_n_396, mul_22_25_n_397, mul_22_25_n_398,
     mul_22_25_n_399, mul_22_25_n_400, mul_22_25_n_401, mul_22_25_n_402,
     mul_22_25_n_403, mul_22_25_n_404, mul_22_25_n_405, mul_22_25_n_406,
     mul_22_25_n_407, mul_22_25_n_408, mul_22_25_n_409, mul_22_25_n_410,
     mul_22_25_n_411, mul_22_25_n_412, mul_22_25_n_413, mul_22_25_n_414,
     mul_22_25_n_415, mul_22_25_n_416, mul_22_25_n_417, mul_22_25_n_418,
     mul_22_25_n_419, mul_22_25_n_420, mul_22_25_n_421, mul_22_25_n_422,
     mul_22_25_n_423, mul_22_25_n_424, mul_22_25_n_425, mul_22_25_n_426,
     mul_22_25_n_427, mul_22_25_n_428, mul_22_25_n_429, mul_22_25_n_430,
     mul_22_25_n_431, mul_22_25_n_432, mul_22_25_n_433, mul_22_25_n_434,
     mul_22_25_n_435, mul_22_25_n_436, mul_22_25_n_437, mul_22_25_n_438,
     mul_22_25_n_439, mul_22_25_n_440, mul_22_25_n_441, mul_22_25_n_442,
     mul_22_25_n_443, mul_22_25_n_444, mul_22_25_n_445, mul_22_25_n_446,
     mul_22_25_n_447, mul_22_25_n_448, mul_22_25_n_449, mul_22_25_n_450,
     mul_22_25_n_451, mul_22_25_n_452, mul_22_25_n_453, mul_22_25_n_454,
     mul_22_25_n_455, mul_22_25_n_456, mul_22_25_n_457, mul_22_25_n_459,
     mul_22_25_n_460, mul_22_25_n_461, mul_22_25_n_462, mul_22_25_n_463,
     mul_22_25_n_464, mul_22_25_n_465, mul_22_25_n_466, mul_22_25_n_467,
     mul_22_25_n_468, mul_22_25_n_469, mul_22_25_n_470, mul_22_25_n_471,
     mul_22_25_n_472, mul_22_25_n_473, mul_22_25_n_474, mul_22_25_n_475,
     mul_22_25_n_476, mul_22_25_n_477, mul_22_25_n_478, mul_22_25_n_479,
     mul_22_25_n_480, mul_22_25_n_481, mul_22_25_n_482, mul_22_25_n_483,
     mul_22_25_n_484, mul_22_25_n_485, mul_22_25_n_486, mul_22_25_n_487,
     mul_22_25_n_488, mul_22_25_n_489, mul_22_25_n_490, mul_22_25_n_491,
     mul_22_25_n_492, mul_22_25_n_493, mul_22_25_n_494, mul_22_25_n_495,
     mul_22_25_n_496, mul_22_25_n_497, mul_22_25_n_498, mul_22_25_n_499,
     mul_22_25_n_500, mul_22_25_n_501, mul_22_25_n_502, mul_22_25_n_503,
     mul_22_25_n_504, mul_22_25_n_505, mul_22_25_n_506, mul_22_25_n_507,
     mul_22_25_n_508, mul_22_25_n_509, mul_22_25_n_510, mul_22_25_n_511,
     mul_22_25_n_512, mul_22_25_n_513, mul_22_25_n_514, mul_22_25_n_515,
     mul_22_25_n_516, mul_22_25_n_517, mul_22_25_n_518, mul_22_25_n_519,
     mul_22_25_n_520, mul_22_25_n_521, mul_22_25_n_522, mul_22_25_n_523,
     mul_22_25_n_524, mul_22_25_n_525, mul_22_25_n_526, mul_22_25_n_527,
     mul_22_25_n_528, mul_22_25_n_529, mul_22_25_n_530, mul_22_25_n_531,
     mul_22_25_n_532, mul_22_25_n_533, mul_22_25_n_534, mul_22_25_n_535,
     mul_22_25_n_536, mul_22_25_n_537, mul_22_25_n_538, mul_22_25_n_539,
     mul_22_25_n_540, mul_22_25_n_541, mul_22_25_n_542, mul_22_25_n_543,
     mul_22_25_n_544, mul_22_25_n_545, mul_22_25_n_546, mul_22_25_n_547,
     mul_22_25_n_548, mul_22_25_n_549, mul_22_25_n_550, mul_22_25_n_551,
     mul_22_25_n_552, mul_22_25_n_553, mul_22_25_n_554, mul_22_25_n_555,
     mul_22_25_n_556, mul_22_25_n_557, mul_22_25_n_558, mul_22_25_n_559,
     mul_22_25_n_560, mul_22_25_n_561, mul_22_25_n_562, mul_22_25_n_563,
     mul_22_25_n_564, mul_22_25_n_565, mul_22_25_n_566, mul_22_25_n_567,
     mul_22_25_n_568, mul_22_25_n_569, mul_22_25_n_570, mul_22_25_n_571,
     mul_22_25_n_572, mul_22_25_n_573, mul_22_25_n_574, mul_22_25_n_575,
     mul_22_25_n_576, mul_22_25_n_577, mul_22_25_n_578, mul_22_25_n_579,
     mul_22_25_n_580, mul_22_25_n_581, mul_22_25_n_582, mul_22_25_n_583,
     mul_22_25_n_584, mul_22_25_n_585, mul_22_25_n_586, mul_22_25_n_587,
     mul_22_25_n_588, mul_22_25_n_589, mul_22_25_n_590, mul_22_25_n_591,
     mul_22_25_n_592, mul_22_25_n_593, mul_22_25_n_594, mul_22_25_n_595,
     mul_22_25_n_596, mul_22_25_n_597, mul_22_25_n_598, mul_22_25_n_599,
     mul_22_25_n_600, mul_22_25_n_601, mul_22_25_n_602, mul_22_25_n_603,
     mul_22_25_n_604, mul_22_25_n_605, mul_22_25_n_606, mul_22_25_n_607,
     mul_22_25_n_608, mul_22_25_n_609, mul_22_25_n_610, mul_22_25_n_611,
     mul_22_25_n_612, mul_22_25_n_613, mul_22_25_n_614, mul_22_25_n_615,
     mul_22_25_n_616, mul_22_25_n_617, mul_22_25_n_618, mul_22_25_n_619,
     mul_22_25_n_620, mul_22_25_n_621, mul_22_25_n_622, mul_22_25_n_623,
     mul_22_25_n_624, mul_22_25_n_625, mul_22_25_n_626, mul_22_25_n_627,
     mul_22_25_n_628, mul_22_25_n_629, mul_22_25_n_630, mul_22_25_n_631,
     mul_22_25_n_632, mul_22_25_n_633, mul_22_25_n_634, mul_22_25_n_635,
     mul_22_25_n_636, mul_22_25_n_637, mul_22_25_n_638, mul_22_25_n_639,
     mul_22_25_n_640, mul_22_25_n_641, mul_22_25_n_642, mul_22_25_n_643,
     mul_22_25_n_644, mul_22_25_n_645, mul_22_25_n_646, mul_22_25_n_647,
     mul_22_25_n_648, mul_22_25_n_649, mul_22_25_n_650, mul_22_25_n_651,
     mul_22_25_n_652, mul_22_25_n_653, mul_22_25_n_654, mul_22_25_n_655,
     mul_22_25_n_656, mul_22_25_n_657, mul_22_25_n_658, mul_22_25_n_659,
     mul_22_25_n_660, mul_22_25_n_661, mul_22_25_n_662, mul_22_25_n_663,
     mul_22_25_n_664, mul_22_25_n_665, mul_22_25_n_666, mul_22_25_n_667,
     mul_22_25_n_668, mul_22_25_n_669, mul_22_25_n_670, mul_22_25_n_671,
     mul_22_25_n_672, mul_22_25_n_673, mul_22_25_n_674, mul_22_25_n_675,
     mul_22_25_n_676, mul_22_25_n_677, mul_22_25_n_678, mul_22_25_n_679,
     mul_22_25_n_680, mul_22_25_n_681, mul_22_25_n_682, mul_22_25_n_683,
     mul_22_25_n_684, mul_22_25_n_685, mul_22_25_n_686, mul_22_25_n_687,
     mul_22_25_n_688, mul_22_25_n_689, mul_22_25_n_690, mul_22_25_n_691,
     mul_22_25_n_692, mul_22_25_n_693, mul_22_25_n_694, mul_22_25_n_695,
     mul_22_25_n_696, mul_22_25_n_697, mul_22_25_n_698, mul_22_25_n_699,
     mul_22_25_n_700, mul_22_25_n_701, mul_22_25_n_702, mul_22_25_n_703,
     mul_22_25_n_704, mul_22_25_n_705, mul_22_25_n_706, mul_22_25_n_707,
     mul_22_25_n_708, mul_22_25_n_709, mul_22_25_n_710, mul_22_25_n_711,
     mul_22_25_n_712, mul_22_25_n_713, mul_22_25_n_714, mul_22_25_n_715,
     mul_22_25_n_716, mul_22_25_n_717, mul_22_25_n_718, mul_22_25_n_719,
     mul_22_25_n_720, mul_22_25_n_721, mul_22_25_n_722, mul_22_25_n_723,
     mul_22_25_n_724, mul_22_25_n_725, mul_22_25_n_726, mul_22_25_n_727,
     mul_22_25_n_728, mul_22_25_n_729, mul_22_25_n_730, mul_22_25_n_731,
     mul_22_25_n_732, mul_22_25_n_733, mul_22_25_n_734, mul_22_25_n_735,
     mul_22_25_n_736, mul_22_25_n_737, mul_22_25_n_738, mul_22_25_n_739,
     mul_22_25_n_740, mul_22_25_n_741, mul_22_25_n_742, mul_22_25_n_743,
     mul_22_25_n_744, mul_22_25_n_745, mul_22_25_n_746, mul_22_25_n_747,
     mul_22_25_n_748, mul_22_25_n_749, mul_22_25_n_750, mul_22_25_n_751,
     mul_22_25_n_752, mul_22_25_n_753, mul_22_25_n_754, mul_22_25_n_755,
     mul_22_25_n_756, mul_22_25_n_757, mul_22_25_n_758, mul_22_25_n_759,
     mul_22_25_n_760, mul_22_25_n_761, mul_22_25_n_762, mul_22_25_n_763,
     mul_22_25_n_764, mul_22_25_n_765, mul_22_25_n_766, mul_22_25_n_767,
     mul_22_25_n_768, mul_22_25_n_769, mul_22_25_n_770, mul_22_25_n_771,
     mul_22_25_n_772, mul_22_25_n_773, mul_22_25_n_774, mul_22_25_n_775,
     mul_22_25_n_776, mul_22_25_n_777, mul_22_25_n_778, mul_22_25_n_779,
     mul_22_25_n_780, mul_22_25_n_781, mul_22_25_n_782, mul_22_25_n_783,
     mul_22_25_n_784, mul_22_25_n_785, mul_22_25_n_786, mul_22_25_n_787,
     mul_22_25_n_788, mul_22_25_n_789, mul_22_25_n_790, mul_22_25_n_791,
     mul_22_25_n_792, mul_22_25_n_793, mul_22_25_n_794, mul_22_25_n_795,
     mul_22_25_n_796, mul_22_25_n_797, mul_22_25_n_798, mul_22_25_n_799,
     mul_22_25_n_800, mul_22_25_n_801, mul_22_25_n_802, mul_22_25_n_803,
     mul_22_25_n_804, mul_22_25_n_805, mul_22_25_n_806, mul_22_25_n_807,
     mul_22_25_n_808, mul_22_25_n_809, mul_22_25_n_810, mul_22_25_n_811,
     mul_22_25_n_812, mul_22_25_n_813, mul_22_25_n_814, mul_22_25_n_815,
     mul_22_25_n_816, mul_22_25_n_817, mul_22_25_n_818, mul_22_25_n_819,
     mul_22_25_n_820, mul_22_25_n_821, mul_22_25_n_822, mul_22_25_n_823,
     mul_22_25_n_824, mul_22_25_n_825, mul_22_25_n_826, mul_22_25_n_827,
     mul_22_25_n_828, mul_22_25_n_829, mul_22_25_n_830, mul_22_25_n_831,
     mul_22_25_n_832, mul_22_25_n_833, mul_22_25_n_834, mul_22_25_n_835,
     mul_22_25_n_836, mul_22_25_n_837, mul_22_25_n_838, mul_22_25_n_839,
     mul_22_25_n_840, mul_22_25_n_841, mul_22_25_n_842, mul_22_25_n_844,
     mul_22_25_n_845, mul_22_25_n_846, mul_22_25_n_847, mul_22_25_n_848,
     mul_22_25_n_849, mul_22_25_n_850, mul_22_25_n_851, mul_22_25_n_852,
     mul_22_25_n_853, mul_22_25_n_854, mul_22_25_n_855, mul_22_25_n_856,
     mul_22_25_n_857, mul_22_25_n_858, mul_22_25_n_859, mul_22_25_n_860,
     mul_22_25_n_861, mul_22_25_n_862, mul_22_25_n_863, mul_22_25_n_864,
     mul_22_25_n_865, mul_22_25_n_866, mul_22_25_n_868, mul_22_25_n_869,
     mul_22_25_n_870, mul_22_25_n_871, mul_22_25_n_872, mul_22_25_n_873,
     mul_22_25_n_874, mul_22_25_n_875, mul_22_25_n_876, mul_22_25_n_877,
     mul_22_25_n_878, mul_22_25_n_879, mul_22_25_n_880, mul_22_25_n_881,
     mul_22_25_n_882, mul_22_25_n_883, mul_22_25_n_884, mul_22_25_n_885,
     mul_22_25_n_886, mul_22_25_n_887, mul_22_25_n_888, mul_22_25_n_889,
     mul_22_25_n_890, mul_22_25_n_891, mul_22_25_n_892, mul_22_25_n_893,
     mul_22_25_n_894, mul_22_25_n_895, mul_22_25_n_896, mul_22_25_n_897,
     mul_22_25_n_898, mul_22_25_n_899, mul_22_25_n_900, mul_22_25_n_901,
     mul_22_25_n_902, mul_22_25_n_903, mul_22_25_n_904, mul_22_25_n_905,
     mul_22_25_n_906, mul_22_25_n_907, mul_22_25_n_908, mul_22_25_n_909,
     mul_22_25_n_910, mul_22_25_n_911, mul_22_25_n_913, mul_22_25_n_914,
     mul_22_25_n_915, mul_22_25_n_916, mul_22_25_n_917, mul_22_25_n_919,
     mul_22_25_n_920, mul_22_25_n_921, mul_22_25_n_922, mul_22_25_n_923,
     mul_22_25_n_924, mul_22_25_n_926, mul_22_25_n_927, mul_22_25_n_928,
     mul_22_25_n_929, mul_22_25_n_930, mul_22_25_n_932, mul_22_25_n_933,
     mul_22_25_n_934, mul_22_25_n_935, mul_22_25_n_936, mul_22_25_n_937,
     mul_22_25_n_938, mul_22_25_n_939, mul_22_25_n_940, mul_22_25_n_941,
     mul_22_25_n_942, mul_22_25_n_943, mul_22_25_n_944, mul_22_25_n_946,
     mul_22_25_n_947, mul_22_25_n_949, mul_22_25_n_950, mul_22_25_n_951,
     mul_22_25_n_952, mul_22_25_n_953, mul_22_25_n_954, mul_22_25_n_955,
     mul_22_25_n_957, mul_22_25_n_958, mul_22_25_n_959, mul_22_25_n_960,
     mul_22_25_n_961, mul_22_25_n_962, mul_22_25_n_963, mul_22_25_n_964,
     mul_22_25_n_965, mul_22_25_n_966, mul_22_25_n_967, mul_22_25_n_968,
     mul_22_25_n_969, mul_22_25_n_970, mul_22_25_n_971, mul_22_25_n_972,
     mul_22_25_n_973, mul_22_25_n_974, mul_22_25_n_975, mul_22_25_n_976,
     mul_22_25_n_977, mul_22_25_n_978, mul_22_25_n_979, mul_22_25_n_980,
     mul_22_25_n_982, mul_22_25_n_983, mul_22_25_n_984, mul_22_25_n_985,
     mul_22_25_n_986, mul_22_25_n_987, mul_22_25_n_988, mul_22_25_n_989,
     mul_22_25_n_990, mul_22_25_n_991, mul_22_25_n_992, mul_22_25_n_993,
     mul_22_25_n_994, mul_22_25_n_995, mul_22_25_n_996, mul_22_25_n_997,
     mul_22_25_n_998, mul_22_25_n_999, mul_22_25_n_1002, mul_22_25_n_1003,
     mul_22_25_n_1004, mul_22_25_n_1005, mul_22_25_n_1006, mul_22_25_n_1007,
     mul_22_25_n_1008, mul_22_25_n_1009, mul_22_25_n_1010, mul_22_25_n_1011,
     mul_22_25_n_1012, mul_22_25_n_1013, mul_22_25_n_1014, mul_22_25_n_1015,
     mul_22_25_n_1016, mul_22_25_n_1017, mul_22_25_n_1018, mul_22_25_n_1019,
     mul_22_25_n_1020, mul_22_25_n_1021, mul_22_25_n_1022, mul_22_25_n_1023,
     mul_22_25_n_1024, mul_22_25_n_1025, mul_22_25_n_1026, mul_22_25_n_1027,
     mul_22_25_n_1028, mul_22_25_n_1029, mul_22_25_n_1030, mul_22_25_n_1031,
     mul_22_25_n_1032, mul_22_25_n_1033, mul_22_25_n_1034, mul_22_25_n_1035,
     mul_22_25_n_1036, mul_22_25_n_1037, mul_22_25_n_1038, mul_22_25_n_1039,
     mul_22_25_n_1040, mul_22_25_n_1041, mul_22_25_n_1042, mul_22_25_n_1044,
     mul_22_25_n_1045, mul_22_25_n_1046, mul_22_25_n_1047, mul_22_25_n_1048,
     mul_22_25_n_1049, mul_22_25_n_1050, mul_22_25_n_1052, mul_22_25_n_1053,
     mul_22_25_n_1054, mul_22_25_n_1055, mul_22_25_n_1056, mul_22_25_n_1057,
     mul_22_25_n_1058, mul_22_25_n_1059, mul_22_25_n_1060, mul_22_25_n_1061,
     mul_22_25_n_1062, mul_22_25_n_1063, mul_22_25_n_1064, mul_22_25_n_1065,
     mul_22_25_n_1066, mul_22_25_n_1067, mul_22_25_n_1068, mul_22_25_n_1069,
     mul_22_25_n_1070, mul_22_25_n_1071, mul_22_25_n_1072, mul_22_25_n_1073,
     mul_22_25_n_1074, mul_22_25_n_1075, mul_22_25_n_1076, mul_22_25_n_1077,
     mul_22_25_n_1078, mul_22_25_n_1079, mul_22_25_n_1080, mul_22_25_n_1081,
     mul_22_25_n_1082, mul_22_25_n_1083, mul_22_25_n_1084, mul_22_25_n_1085,
     mul_22_25_n_1087, mul_22_25_n_1088, mul_22_25_n_1089, mul_22_25_n_1090,
     mul_22_25_n_1091, mul_22_25_n_1092, mul_22_25_n_1093, mul_22_25_n_1094,
     mul_22_25_n_1095, mul_22_25_n_1096, mul_22_25_n_1097, mul_22_25_n_1098,
     mul_22_25_n_1099, mul_22_25_n_1100, mul_22_25_n_1101, mul_22_25_n_1102,
     mul_22_25_n_1103, mul_22_25_n_1104, mul_22_25_n_1105, mul_22_25_n_1106,
     mul_22_25_n_1107, mul_22_25_n_1108, mul_22_25_n_1109, mul_22_25_n_1110,
     mul_22_25_n_1111, mul_22_25_n_1112, mul_22_25_n_1113, mul_22_25_n_1114,
     mul_22_25_n_1115, mul_22_25_n_1116, mul_22_25_n_1117, mul_22_25_n_1118,
     mul_22_25_n_1119, mul_22_25_n_1120, mul_22_25_n_1121, mul_22_25_n_1122,
     mul_22_25_n_1123, mul_22_25_n_1124, mul_22_25_n_1125, mul_22_25_n_1126,
     mul_22_25_n_1127, mul_22_25_n_1128, mul_22_25_n_1129, mul_22_25_n_1130,
     mul_22_25_n_1131, mul_22_25_n_1132, mul_22_25_n_1133, mul_22_25_n_1134,
     mul_22_25_n_1135, mul_22_25_n_1136, mul_22_25_n_1137, mul_22_25_n_1138,
     mul_22_25_n_1139, mul_22_25_n_1140, mul_22_25_n_1142, mul_22_25_n_1143,
     mul_22_25_n_1144, mul_22_25_n_1145, mul_22_25_n_1146, mul_22_25_n_1147,
     mul_22_25_n_1148, mul_22_25_n_1149, mul_22_25_n_1150, mul_22_25_n_1151,
     mul_22_25_n_1152, mul_22_25_n_1153, mul_22_25_n_1154, mul_22_25_n_1155,
     mul_22_25_n_1156, mul_22_25_n_1157, mul_22_25_n_1158, mul_22_25_n_1159,
     mul_22_25_n_1160, mul_22_25_n_1161, mul_22_25_n_1162, mul_22_25_n_1163,
     mul_22_25_n_1164, mul_22_25_n_1165, mul_22_25_n_1166, mul_22_25_n_1167,
     mul_22_25_n_1168, mul_22_25_n_1169, mul_22_25_n_1170, mul_22_25_n_1171,
     mul_22_25_n_1172, mul_22_25_n_1173, mul_22_25_n_1174, mul_22_25_n_1175,
     mul_22_25_n_1176, mul_22_25_n_1177, mul_22_25_n_1178, mul_22_25_n_1179,
     mul_22_25_n_1180, mul_22_25_n_1182, mul_22_25_n_1183, mul_22_25_n_1184,
     mul_22_25_n_1185, mul_22_25_n_1186, mul_22_25_n_1187, mul_22_25_n_1188,
     mul_22_25_n_1189, mul_22_25_n_1190, mul_22_25_n_1191, mul_22_25_n_1192,
     mul_22_25_n_1193, mul_22_25_n_1194, mul_22_25_n_1195, mul_22_25_n_1196,
     mul_22_25_n_1198, mul_22_25_n_1200, mul_22_25_n_1201, mul_22_25_n_1202,
     mul_22_25_n_1203, mul_22_25_n_1204, mul_22_25_n_1205, mul_22_25_n_1206,
     mul_22_25_n_1210, mul_22_25_n_1211, mul_22_25_n_1212, mul_22_25_n_1213,
     mul_22_25_n_1214, mul_22_25_n_1215, mul_22_25_n_1216, mul_22_25_n_1217,
     mul_22_25_n_1218, mul_22_25_n_1224, mul_22_25_n_1225, mul_22_25_n_1226,
     mul_22_25_n_1227, mul_22_25_n_1228, mul_22_25_n_1229, mul_22_25_n_1230,
     mul_22_25_n_1231, mul_22_25_n_1232, mul_22_25_n_1233, mul_22_25_n_1240,
     mul_22_25_n_1241, mul_22_25_n_1242, mul_22_25_n_1243, mul_22_25_n_1245,
     mul_22_25_n_1246, mul_22_25_n_1247, mul_22_25_n_1254, mul_22_25_n_1255,
     mul_22_25_n_1257, mul_22_25_n_1263, mul_22_25_n_1265, mul_22_25_n_1266,
     mul_22_25_n_1267, mul_22_25_n_1268, mul_22_25_n_1269, mul_22_25_n_1270,
     mul_22_25_n_1271, mul_22_25_n_1272, mul_22_25_n_1273, mul_22_25_n_1274,
     mul_22_25_n_1275, mul_22_25_n_1276, mul_22_25_n_1277, mul_22_25_n_1278,
     mul_22_25_n_1279, mul_22_25_n_1280, mul_22_25_n_1281, mul_22_25_n_1282,
     mul_22_25_n_1283, mul_22_25_n_1284, mul_22_25_n_1285, mul_22_25_n_1286,
     mul_22_25_n_1287, mul_22_25_n_1288, mul_22_25_n_1289, mul_22_25_n_1290,
     mul_22_25_n_1291, mul_22_25_n_1292, mul_22_25_n_1293, mul_22_25_n_1294,
     mul_22_25_n_1295, mul_22_25_n_1296, mul_22_25_n_1297, mul_22_25_n_1298,
     mul_22_25_n_1299, mul_22_25_n_1300, mul_22_25_n_1301, mul_22_25_n_1302,
     mul_22_25_n_1303, mul_22_25_n_1304, mul_22_25_n_1305, mul_22_25_n_1306,
     mul_22_25_n_1307, mul_22_25_n_1308, mul_22_25_n_1309, mul_22_25_n_1310,
     mul_22_25_n_1311, mul_22_25_n_1312, mul_22_25_n_1313, mul_22_25_n_1314,
     mul_22_25_n_1315, mul_22_25_n_1316, mul_22_25_n_1317, mul_22_25_n_1318,
     mul_22_25_n_1319, mul_22_25_n_1320, mul_22_25_n_1321, mul_22_25_n_1322,
     mul_22_25_n_1323, mul_22_25_n_1324, mul_22_25_n_1325, mul_22_25_n_1326,
     mul_22_25_n_1327, mul_22_25_n_1328, mul_22_25_n_1329, mul_22_25_n_1330,
     mul_22_25_n_1331, mul_22_25_n_1332, mul_22_25_n_1333, mul_22_25_n_1334,
     mul_22_25_n_1335, mul_22_25_n_1336, mul_22_25_n_1337, mul_22_25_n_1338,
     mul_22_25_n_1339, mul_22_25_n_1340, mul_22_25_n_1341, mul_22_25_n_1342,
     mul_22_25_n_1343, mul_22_25_n_1344, mul_22_25_n_1345, mul_22_25_n_1346,
     mul_22_25_n_1347, mul_22_25_n_1348, mul_22_25_n_1349, mul_22_25_n_1350,
     mul_22_25_n_1351, mul_22_25_n_1352, mul_22_25_n_1353, mul_22_25_n_1354,
     mul_22_25_n_1355, mul_22_25_n_1356, mul_22_25_n_1357, mul_22_25_n_1358,
     mul_22_25_n_1359, mul_22_25_n_1360, mul_22_25_n_1361, mul_22_25_n_1362,
     mul_22_25_n_1363, mul_22_25_n_1364, mul_22_25_n_1365, mul_22_25_n_1366,
     mul_22_25_n_1367, mul_22_25_n_1368, mul_22_25_n_1369, mul_22_25_n_1370,
     mul_22_25_n_1371, mul_22_25_n_1372, mul_22_25_n_1373, mul_22_25_n_1374,
     mul_22_25_n_1375, mul_22_25_n_1376, mul_22_25_n_1377, mul_22_25_n_1378,
     mul_22_25_n_1379, mul_22_25_n_1380, mul_22_25_n_1381, mul_22_25_n_1382,
     mul_22_25_n_1383, mul_22_25_n_1384, mul_22_25_n_1385, mul_22_25_n_1386,
     mul_22_25_n_1387, mul_22_25_n_1388, mul_22_25_n_1389, mul_22_25_n_1390,
     mul_22_25_n_1391, mul_22_25_n_1392, mul_22_25_n_1393, mul_22_25_n_1394,
     mul_22_25_n_1395, mul_22_25_n_1396, mul_22_25_n_1397, mul_22_25_n_1398,
     mul_22_25_n_1399, mul_22_25_n_1400, mul_22_25_n_1401, mul_22_25_n_1402,
     mul_22_25_n_1403, mul_22_25_n_1404, mul_22_25_n_1405, mul_22_25_n_1406,
     mul_22_25_n_1407, mul_22_25_n_1408, mul_22_25_n_1409, mul_22_25_n_1410,
     mul_22_25_n_1411, mul_22_25_n_1412, mul_22_25_n_1413, mul_22_25_n_1414,
     mul_22_25_n_1415, mul_22_25_n_1416, mul_22_25_n_1417, mul_22_25_n_1418,
     mul_22_25_n_1419, mul_22_25_n_1420, mul_22_25_n_1421, mul_22_25_n_1422,
     mul_22_25_n_1423, mul_22_25_n_1424, mul_22_25_n_1425, mul_22_25_n_1426,
     mul_22_25_n_1427, mul_22_25_n_1428, mul_22_25_n_1429, mul_22_25_n_1430,
     mul_22_25_n_1431, mul_22_25_n_1432, mul_22_25_n_1433, mul_22_25_n_1434,
     mul_22_25_n_1435, mul_22_25_n_1436, mul_22_25_n_1437, mul_22_25_n_1438,
     mul_22_25_n_1439, mul_22_25_n_1440, mul_22_25_n_1441, mul_22_25_n_1442,
     mul_22_25_n_1443, mul_22_25_n_1444, mul_22_25_n_1445, mul_22_25_n_1446,
     mul_22_25_n_1447, mul_22_25_n_1448, mul_22_25_n_1449, mul_22_25_n_1450,
     mul_22_25_n_1451, mul_22_25_n_1452, mul_22_25_n_1453, mul_22_25_n_1454,
     mul_22_25_n_1455, mul_22_25_n_1456, mul_22_25_n_1457, mul_22_25_n_1458,
     mul_22_25_n_1459, mul_22_25_n_1460, mul_22_25_n_1461, mul_22_25_n_1462,
     mul_22_25_n_1463, mul_22_25_n_1464, mul_22_25_n_1465, mul_22_25_n_1466,
     mul_22_25_n_1467, mul_22_25_n_1468, mul_22_25_n_1469, mul_22_25_n_1470,
     mul_22_25_n_1471, mul_22_25_n_1472, mul_22_25_n_1473, mul_22_25_n_1474,
     mul_22_25_n_1475, mul_22_25_n_1476, mul_22_25_n_1477, mul_22_25_n_1478,
     mul_22_25_n_1479, mul_22_25_n_1480, mul_22_25_n_1481, mul_22_25_n_1482,
     mul_22_25_n_1483, mul_22_25_n_1484, mul_22_25_n_1485, mul_22_25_n_1486,
     mul_22_25_n_1487, mul_22_25_n_1488, mul_22_25_n_1489, mul_22_25_n_1490,
     mul_22_25_n_1491, mul_22_25_n_1492, mul_22_25_n_1493, mul_22_25_n_1494,
     mul_22_25_n_1495, mul_22_25_n_1496, mul_22_25_n_1497, mul_22_25_n_1498,
     mul_22_25_n_1499, mul_22_25_n_1500, mul_22_25_n_1501, mul_22_25_n_1502,
     mul_22_25_n_1503, mul_22_25_n_1504, mul_22_25_n_1505, mul_22_25_n_1506,
     mul_22_25_n_1507, mul_22_25_n_1508, mul_22_25_n_1509, mul_22_25_n_1510,
     mul_22_25_n_1511, mul_22_25_n_1512, mul_22_25_n_1513, mul_22_25_n_1514,
     mul_22_25_n_1515, mul_22_25_n_1516, mul_22_25_n_1517, mul_22_25_n_1518,
     mul_22_25_n_1519, mul_22_25_n_1520, mul_22_25_n_1521, mul_22_25_n_1522,
     mul_22_25_n_1523, mul_22_25_n_1524, mul_22_25_n_1525, mul_22_25_n_1526,
     mul_22_25_n_1527, mul_22_25_n_1528, mul_22_25_n_1529, mul_22_25_n_1530,
     mul_22_25_n_1531, mul_22_25_n_1532, mul_22_25_n_1533, mul_22_25_n_1534,
     mul_22_25_n_1535, mul_22_25_n_1536, mul_22_25_n_1537, mul_22_25_n_1538,
     mul_22_25_n_1539, mul_22_25_n_1540, mul_22_25_n_1541, mul_22_25_n_1542,
     mul_22_25_n_1543, mul_22_25_n_1544, mul_22_25_n_1545, mul_22_25_n_1546,
     mul_22_25_n_1547, mul_22_25_n_1548, mul_22_25_n_1549, mul_22_25_n_1550,
     mul_22_25_n_1551, mul_22_25_n_1552, mul_22_25_n_1553, mul_22_25_n_1554,
     mul_22_25_n_1555, mul_22_25_n_1556, mul_22_25_n_1557, mul_22_25_n_1558,
     mul_22_25_n_1559, mul_22_25_n_1560, mul_22_25_n_1561, mul_22_25_n_1562,
     mul_22_25_n_1563, mul_22_25_n_1564, mul_22_25_n_1565, mul_22_25_n_1566,
     mul_22_25_n_1567, mul_22_25_n_1568, mul_22_25_n_1569, mul_22_25_n_1570,
     mul_22_25_n_1571, mul_22_25_n_1572, mul_22_25_n_1573, mul_22_25_n_1574,
     mul_22_25_n_1575, mul_22_25_n_1576, mul_22_25_n_1577, mul_22_25_n_1578,
     mul_22_25_n_1579, mul_22_25_n_1580, mul_22_25_n_1581, mul_22_25_n_1582,
     mul_22_25_n_1583, mul_22_25_n_1584, mul_22_25_n_1585, mul_22_25_n_1586,
     mul_22_25_n_1587, mul_22_25_n_1588, mul_22_25_n_1589, mul_22_25_n_1590,
     mul_22_25_n_1591, mul_22_25_n_1592, mul_22_25_n_1593, mul_22_25_n_1594,
     mul_22_25_n_1595, mul_22_25_n_1596, mul_22_25_n_1597, mul_22_25_n_1598,
     mul_22_25_n_1599, mul_22_25_n_1600, mul_22_25_n_1601, mul_22_25_n_1602,
     mul_22_25_n_1603, mul_22_25_n_1604, mul_22_25_n_1605, mul_22_25_n_1606,
     mul_22_25_n_1607, mul_22_25_n_1608, mul_22_25_n_1609, mul_22_25_n_1610,
     mul_22_25_n_1611, mul_22_25_n_1612, mul_22_25_n_1613, mul_22_25_n_1614,
     mul_22_25_n_1615, mul_22_25_n_1616, mul_22_25_n_1617, mul_22_25_n_1618,
     mul_22_25_n_1619, mul_22_25_n_1620, mul_22_25_n_1621, mul_22_25_n_1622,
     mul_22_25_n_1623, mul_22_25_n_1624, mul_22_25_n_1625, mul_22_25_n_1626,
     mul_22_25_n_1627, mul_22_25_n_1628, mul_22_25_n_1629, mul_22_25_n_1630,
     mul_22_25_n_1631, mul_22_25_n_1632, mul_22_25_n_1633, mul_22_25_n_1634,
     mul_22_25_n_1635, mul_22_25_n_1636, mul_22_25_n_1637, mul_22_25_n_1638,
     mul_22_25_n_1639, mul_22_25_n_1640, mul_22_25_n_1641, mul_22_25_n_1642,
     mul_22_25_n_1643, mul_22_25_n_1644, mul_22_25_n_1645, mul_22_25_n_1646,
     mul_22_25_n_1647, mul_22_25_n_1648, mul_22_25_n_1649, mul_22_25_n_1650,
     mul_22_25_n_1651, mul_22_25_n_1652, mul_22_25_n_1653, mul_22_25_n_1654,
     mul_22_25_n_1655, mul_22_25_n_1656, mul_22_25_n_1657, mul_22_25_n_1658,
     mul_22_25_n_1659, mul_22_25_n_1660, mul_22_25_n_1661, mul_22_25_n_1662,
     mul_22_25_n_1663, mul_22_25_n_1664, mul_22_25_n_1665, mul_22_25_n_1666,
     mul_22_25_n_1667, mul_22_25_n_1668, mul_22_25_n_1669, mul_22_25_n_1670,
     mul_22_25_n_1671, mul_22_25_n_1672, mul_22_25_n_1673, mul_22_25_n_1674,
     mul_22_25_n_1675, mul_22_25_n_1676, mul_22_25_n_1677, mul_22_25_n_1678,
     mul_22_25_n_1679, mul_22_25_n_1680, mul_22_25_n_1681, mul_22_25_n_1682,
     mul_22_25_n_1683, mul_22_25_n_1684, mul_22_25_n_1685, mul_22_25_n_1686,
     mul_22_25_n_1687, mul_22_25_n_1688, mul_22_25_n_1689, mul_22_25_n_1690,
     mul_22_25_n_1691, mul_22_25_n_1692, mul_22_25_n_1693, mul_22_25_n_1694,
     mul_22_25_n_1695, mul_22_25_n_1696, mul_22_25_n_1697, mul_22_25_n_1698,
     mul_22_25_n_1699, mul_22_25_n_1700, mul_22_25_n_1701, mul_22_25_n_1702,
     mul_22_25_n_1703, mul_22_25_n_1704, mul_22_25_n_1705, mul_22_25_n_1706,
     mul_22_25_n_1707, mul_22_25_n_1708, mul_22_25_n_1709, mul_22_25_n_1710,
     mul_22_25_n_1711, mul_22_25_n_1712, mul_22_25_n_1713, mul_22_25_n_1714,
     mul_22_25_n_1715, mul_22_25_n_1716, mul_22_25_n_1717, mul_22_25_n_1718,
     mul_22_25_n_1719, mul_22_25_n_1720, mul_22_25_n_1721, mul_22_25_n_1722,
     mul_22_25_n_1723, mul_22_25_n_1724, mul_22_25_n_1725, mul_22_25_n_1726,
     mul_22_25_n_1727, mul_22_25_n_1728, mul_22_25_n_1729, mul_22_25_n_1730,
     mul_22_25_n_1731, mul_22_25_n_1732, mul_22_25_n_1733, mul_22_25_n_1734,
     mul_22_25_n_1735, mul_22_25_n_1736, mul_22_25_n_1737, mul_22_25_n_1738,
     mul_22_25_n_1739, mul_22_25_n_1740, mul_22_25_n_1741, mul_22_25_n_1742,
     mul_22_25_n_1743, mul_22_25_n_1744, mul_22_25_n_1745, mul_22_25_n_1746,
     mul_22_25_n_1747, mul_22_25_n_1748, mul_22_25_n_1749, mul_22_25_n_1750,
     mul_22_25_n_1751, mul_22_25_n_1752, mul_22_25_n_1753, mul_22_25_n_1754,
     mul_22_25_n_1755, mul_22_25_n_1756, mul_22_25_n_1757, mul_22_25_n_1758,
     mul_22_25_n_1759, mul_22_25_n_1760, mul_22_25_n_1761, mul_22_25_n_1762,
     mul_22_25_n_1763, mul_22_25_n_1764, mul_22_25_n_1765, mul_22_25_n_1766,
     mul_22_25_n_1767, mul_22_25_n_1768, mul_22_25_n_1769, mul_22_25_n_1770,
     mul_22_25_n_1771, mul_22_25_n_1772, mul_22_25_n_1773, mul_22_25_n_1774,
     mul_22_25_n_1775, mul_22_25_n_1776, mul_22_25_n_1777, mul_22_25_n_1778,
     mul_22_25_n_1779, mul_22_25_n_1780, mul_22_25_n_1781, mul_22_25_n_1782,
     mul_22_25_n_1783, mul_22_25_n_1784, mul_22_25_n_1785, mul_22_25_n_1786,
     mul_22_25_n_1787, mul_22_25_n_1788, mul_22_25_n_1789, mul_22_25_n_1790,
     mul_22_25_n_1791, mul_22_25_n_1792, mul_22_25_n_1793, mul_22_25_n_1794,
     mul_22_25_n_1795, mul_22_25_n_1796, mul_22_25_n_1797, mul_22_25_n_1798,
     mul_22_25_n_1799, mul_22_25_n_1800, mul_22_25_n_1801, mul_22_25_n_1802,
     mul_22_25_n_1803, mul_22_25_n_1804, mul_22_25_n_1805, mul_22_25_n_1806,
     mul_22_25_n_1807, mul_22_25_n_1808, mul_22_25_n_1809, mul_22_25_n_1810,
     mul_22_25_n_1811, mul_22_25_n_1812, mul_22_25_n_1813, mul_22_25_n_1814,
     mul_22_25_n_1815, mul_22_25_n_1816, mul_22_25_n_1817, mul_22_25_n_1818,
     mul_22_25_n_1819, n_0, n_42, n_43, n_44, n_45, n_46, n_47, n_48, n_51, n_55,
     n_57, n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_68, n_69, n_71, n_72,
     n_73, n_74, n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_84,
     n_85, n_86, n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96,
     n_97, n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107,
     n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118,
     n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129,
     n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140,
     n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151,
     n_152, clk, clr, n_210, asc001_0_, asc001_1_, asc001_2_, asc001_3_,
     asc001_4_, asc001_5_, asc001_6_, asc001_7_, asc001_8_, asc001_9_,
     asc001_10_, asc001_11_, asc001_12_, asc001_13_, asc001_14_, asc001_15_,
     asc001_16_, asc001_17_, asc001_18_, asc001_19_, asc001_20_, asc001_21_,
     asc001_22_, asc001_23_, asc001_24_, asc001_25_, asc001_26_, asc001_27_,
     asc001_28_, asc001_29_, asc001_30_, asc001_31_, asc001_32_, asc001_33_,
     asc001_34_, asc001_35_, asc001_36_, asc001_37_, asc001_38_, asc001_39_,
     asc001_40_, asc001_41_, asc001_42_, asc001_43_, asc001_44_, asc001_45_,
     asc001_46_, asc001_47_, asc001_48_, asc001_49_;
assign {out1[49]} = asc001_49_;
assign {out1[48]} = asc001_48_;
assign {out1[47]} = asc001_47_;
assign {out1[46]} = asc001_46_;
assign {out1[45]} = asc001_45_;
assign {out1[44]} = asc001_44_;
assign {out1[43]} = asc001_43_;
assign {out1[42]} = asc001_42_;
assign {out1[41]} = asc001_41_;
assign {out1[40]} = asc001_40_;
assign {out1[39]} = asc001_39_;
assign {out1[38]} = asc001_38_;
assign {out1[37]} = asc001_37_;
assign {out1[36]} = asc001_36_;
assign {out1[35]} = asc001_35_;
assign {out1[34]} = asc001_34_;
assign {out1[33]} = asc001_33_;
assign {out1[32]} = asc001_32_;
assign {out1[31]} = asc001_31_;
assign {out1[30]} = asc001_30_;
assign {out1[29]} = asc001_29_;
assign {out1[28]} = asc001_28_;
assign {out1[27]} = asc001_27_;
assign {out1[26]} = asc001_26_;
assign {out1[25]} = asc001_25_;
assign {out1[24]} = asc001_24_;
assign {out1[23]} = asc001_23_;
assign {out1[22]} = asc001_22_;
assign {out1[21]} = asc001_21_;
assign {out1[20]} = asc001_20_;
assign {out1[19]} = asc001_19_;
assign {out1[18]} = asc001_18_;
assign {out1[17]} = asc001_17_;
assign {out1[16]} = asc001_16_;
assign {out1[15]} = asc001_15_;
assign {out1[14]} = asc001_14_;
assign {out1[13]} = asc001_13_;
assign {out1[12]} = asc001_12_;
assign {out1[11]} = asc001_11_;
assign {out1[10]} = asc001_10_;
assign {out1[9]} = asc001_9_;
 reg out1_41_L0_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) out1_41_L0_reg_IQ <= 1'B0;
     else begin
         out1_41_L0_reg_IQ <= asc001_8_;
     end
 assign {out1[8]} = out1_41_L0_reg_IQ;
 reg retime_s1_24_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_24_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_24_reg_reg_IQ <= mul_22_25_n_1390;
     end
 assign n_129 = retime_s1_24_reg_reg_IQ;
 reg retime_s1_101_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_101_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_101_reg_reg_IQ <= mul_22_25_n_1014;
     end
 assign n_43 = retime_s1_101_reg_reg_IQ;
 reg retime_s1_26_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_26_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_26_reg_reg_IQ <= mul_22_25_n_1009;
     end
 assign n_127 = retime_s1_26_reg_reg_IQ;
 reg retime_s1_29_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_29_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_29_reg_reg_IQ <= mul_22_25_n_1596;
     end
 assign n_124 = retime_s1_29_reg_reg_IQ;
 reg retime_s1_30_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_30_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_30_reg_reg_IQ <= mul_22_25_n_1613;
     end
 assign n_123 = retime_s1_30_reg_reg_IQ;
 reg retime_s1_34_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_34_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_34_reg_reg_IQ <= mul_22_25_n_1037;
     end
 assign n_119 = retime_s1_34_reg_reg_IQ;
 reg retime_s1_35_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_35_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_35_reg_reg_IQ <= mul_22_25_n_1792;
     end
 assign n_118 = retime_s1_35_reg_reg_IQ;
 reg retime_s1_39_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_39_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_39_reg_reg_IQ <= mul_22_25_n_1012;
     end
 assign n_114 = retime_s1_39_reg_reg_IQ;
 reg retime_s1_40_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_40_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_40_reg_reg_IQ <= mul_22_25_n_1629;
     end
 assign n_113 = retime_s1_40_reg_reg_IQ;
 reg retime_s1_42_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_42_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_42_reg_reg_IQ <= mul_22_25_n_1581;
     end
 assign n_111 = retime_s1_42_reg_reg_IQ;
 reg retime_s1_44_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_44_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_44_reg_reg_IQ <= mul_22_25_n_1002;
     end
 assign n_109 = retime_s1_44_reg_reg_IQ;
 reg retime_s1_47_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_47_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_47_reg_reg_IQ <= mul_22_25_n_1376;
     end
 assign n_106 = retime_s1_47_reg_reg_IQ;
 reg retime_s1_51_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_51_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_51_reg_reg_IQ <= mul_22_25_n_958;
     end
 assign n_102 = retime_s1_51_reg_reg_IQ;
 reg retime_s1_53_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_53_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_53_reg_reg_IQ <= mul_22_25_n_1565;
     end
 assign n_100 = retime_s1_53_reg_reg_IQ;
 reg retime_s1_55_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_55_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_55_reg_reg_IQ <= mul_22_25_n_1549;
     end
 assign n_98 = retime_s1_55_reg_reg_IQ;
 reg retime_s1_57_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_57_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_57_reg_reg_IQ <= mul_22_25_n_1517;
     end
 assign n_96 = retime_s1_57_reg_reg_IQ;
 reg retime_s1_60_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_60_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_60_reg_reg_IQ <= mul_22_25_n_1005;
     end
 assign n_93 = retime_s1_60_reg_reg_IQ;
 reg retime_s1_61_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_61_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_61_reg_reg_IQ <= mul_22_25_n_11;
     end
 assign n_92 = retime_s1_61_reg_reg_IQ;
 reg retime_s1_64_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_64_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_64_reg_reg_IQ <= mul_22_25_n_1405;
     end
 assign n_89 = retime_s1_64_reg_reg_IQ;
 reg retime_s1_75_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_75_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_75_reg_reg_IQ <= mul_22_25_n_983;
     end
 assign n_78 = retime_s1_75_reg_reg_IQ;
 reg retime_s1_77_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_77_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_77_reg_reg_IQ <= mul_22_25_n_1017;
     end
 assign n_76 = retime_s1_77_reg_reg_IQ;
 reg retime_s1_79_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_79_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_79_reg_reg_IQ <= mul_22_25_n_1006;
     end
 assign n_74 = retime_s1_79_reg_reg_IQ;
 reg retime_s1_81_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_81_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_81_reg_reg_IQ <= mul_22_25_n_964;
     end
 assign n_72 = retime_s1_81_reg_reg_IQ;
 reg retime_s1_82_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_82_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_82_reg_reg_IQ <= mul_22_25_n_8;
     end
 assign n_71 = retime_s1_82_reg_reg_IQ;
 reg retime_s1_87_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_87_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_87_reg_reg_IQ <= mul_22_25_n_971;
     end
 assign n_62 = retime_s1_87_reg_reg_IQ;
 reg retime_s1_90_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_90_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_90_reg_reg_IQ <= mul_22_25_n_1453;
     end
 assign n_59 = retime_s1_90_reg_reg_IQ;
 reg retime_s1_95_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_95_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_95_reg_reg_IQ <= mul_22_25_n_1066;
     end
 assign n_51 = retime_s1_95_reg_reg_IQ;
 reg retime_s1_97_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_97_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_97_reg_reg_IQ <= mul_22_25_n_1421;
     end
 assign n_47 = retime_s1_97_reg_reg_IQ;
 reg retime_s1_98_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_98_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_98_reg_reg_IQ <= mul_22_25_n_1437;
     end
 assign n_46 = retime_s1_98_reg_reg_IQ;
 reg retime_s1_100_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_100_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_100_reg_reg_IQ <= mul_22_25_n_965;
     end
 assign n_44 = retime_s1_100_reg_reg_IQ;
 reg retime_s1_102_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_102_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_102_reg_reg_IQ <= mul_22_25_n_1007;
     end
 assign n_42 = retime_s1_102_reg_reg_IQ;
 reg out1_42_L0_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) out1_42_L0_reg_IQ <= 1'B0;
     else begin
         out1_42_L0_reg_IQ <= asc001_7_;
     end
 assign {out1[7]} = out1_42_L0_reg_IQ;
 reg out1_43_L0_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) out1_43_L0_reg_IQ <= 1'B0;
     else begin
         out1_43_L0_reg_IQ <= asc001_6_;
     end
 assign {out1[6]} = out1_43_L0_reg_IQ;
 reg out1_44_L0_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) out1_44_L0_reg_IQ <= 1'B0;
     else begin
         out1_44_L0_reg_IQ <= asc001_5_;
     end
 assign {out1[5]} = out1_44_L0_reg_IQ;
 reg out1_45_L0_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) out1_45_L0_reg_IQ <= 1'B0;
     else begin
         out1_45_L0_reg_IQ <= asc001_4_;
     end
 assign {out1[4]} = out1_45_L0_reg_IQ;
 reg out1_46_L0_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) out1_46_L0_reg_IQ <= 1'B0;
     else begin
         out1_46_L0_reg_IQ <= asc001_3_;
     end
 assign {out1[3]} = out1_46_L0_reg_IQ;
 reg out1_47_L0_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) out1_47_L0_reg_IQ <= 1'B0;
     else begin
         out1_47_L0_reg_IQ <= asc001_2_;
     end
 assign {out1[2]} = out1_47_L0_reg_IQ;
 reg out1_48_L0_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) out1_48_L0_reg_IQ <= 1'B0;
     else begin
         out1_48_L0_reg_IQ <= asc001_1_;
     end
 assign {out1[1]} = out1_48_L0_reg_IQ;
 reg out1_49_L0_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) out1_49_L0_reg_IQ <= 1'B0;
     else begin
         out1_49_L0_reg_IQ <= asc001_0_;
     end
 assign {out1[0]} = out1_49_L0_reg_IQ;
 reg retime_s1_1_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_1_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_1_reg_reg_IQ <= mul_22_25_n_938;
     end
 assign n_152 = retime_s1_1_reg_reg_IQ;
 reg retime_s1_3_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_3_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_3_reg_reg_IQ <= mul_22_25_n_1813;
     end
 assign n_150 = retime_s1_3_reg_reg_IQ;
 reg retime_s1_5_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_5_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_5_reg_reg_IQ <= mul_22_25_n_1363;
     end
 assign n_148 = retime_s1_5_reg_reg_IQ;
 reg retime_s1_6_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_6_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_6_reg_reg_IQ <= mul_22_25_n_1351;
     end
 assign n_147 = retime_s1_6_reg_reg_IQ;
 reg retime_s1_7_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_7_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_7_reg_reg_IQ <= mul_22_25_n_977;
     end
 assign n_146 = retime_s1_7_reg_reg_IQ;
 reg retime_s1_9_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_9_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_9_reg_reg_IQ <= mul_22_25_n_1089;
     end
 assign n_144 = retime_s1_9_reg_reg_IQ;
 reg retime_s1_11_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_11_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_11_reg_reg_IQ <= mul_22_25_n_1501;
     end
 assign n_142 = retime_s1_11_reg_reg_IQ;
 reg retime_s1_13_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_13_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_13_reg_reg_IQ <= mul_22_25_n_1485;
     end
 assign n_140 = retime_s1_13_reg_reg_IQ;
 reg retime_s1_14_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_14_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_14_reg_reg_IQ <= mul_22_25_n_962;
     end
 assign n_139 = retime_s1_14_reg_reg_IQ;
 reg retime_s1_17_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_17_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_17_reg_reg_IQ <= mul_22_25_n_1469;
     end
 assign n_136 = retime_s1_17_reg_reg_IQ;
 reg retime_s1_20_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_20_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_20_reg_reg_IQ <= mul_22_25_n_1533;
     end
 assign n_133 = retime_s1_20_reg_reg_IQ;
 reg retime_s1_23_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_23_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_23_reg_reg_IQ <= mul_22_25_n_1375;
     end
 assign n_130 = retime_s1_23_reg_reg_IQ;
 reg retime_s1_25_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_25_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_25_reg_reg_IQ <= mul_22_25_n_1010;
     end
 assign n_128 = retime_s1_25_reg_reg_IQ;
 reg retime_s1_49_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_49_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_49_reg_reg_IQ <= mul_22_25_n_1377;
     end
 assign n_104 = retime_s1_49_reg_reg_IQ;
 reg retime_s1_18_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_18_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_18_reg_reg_IQ <= mul_22_25_n_1550;
     end
 assign n_135 = retime_s1_18_reg_reg_IQ;
 reg retime_s1_28_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_28_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_28_reg_reg_IQ <= mul_22_25_n_1628;
     end
 assign n_125 = retime_s1_28_reg_reg_IQ;
 reg retime_s1_31_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_31_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_31_reg_reg_IQ <= mul_22_25_n_1580;
     end
 assign n_122 = retime_s1_31_reg_reg_IQ;
 reg retime_s1_32_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_32_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_32_reg_reg_IQ <= mul_22_25_n_1597;
     end
 assign n_121 = retime_s1_32_reg_reg_IQ;
 reg retime_s1_33_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_33_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_33_reg_reg_IQ <= mul_22_25_n_1757;
     end
 assign n_120 = retime_s1_33_reg_reg_IQ;
 reg retime_s1_22_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_22_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_22_reg_reg_IQ <= mul_22_25_n_963;
     end
 assign n_131 = retime_s1_22_reg_reg_IQ;
 reg retime_s1_36_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_36_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_36_reg_reg_IQ <= mul_22_25_n_1470;
     end
 assign n_117 = retime_s1_36_reg_reg_IQ;
 reg retime_s1_37_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_37_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_37_reg_reg_IQ <= mul_22_25_n_1018;
     end
 assign n_116 = retime_s1_37_reg_reg_IQ;
 reg retime_s1_38_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_38_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_38_reg_reg_IQ <= mul_22_25_n_1016;
     end
 assign n_115 = retime_s1_38_reg_reg_IQ;
 reg retime_s1_41_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_41_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_41_reg_reg_IQ <= mul_22_25_n_1564;
     end
 assign n_112 = retime_s1_41_reg_reg_IQ;
 reg retime_s1_96_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_96_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_96_reg_reg_IQ <= mul_22_25_n_1566;
     end
 assign n_48 = retime_s1_96_reg_reg_IQ;
 reg retime_s1_43_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_43_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_43_reg_reg_IQ <= mul_22_25_n_1019;
     end
 assign n_110 = retime_s1_43_reg_reg_IQ;
 reg retime_s1_45_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_45_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_45_reg_reg_IQ <= mul_22_25_n_12;
     end
 assign n_108 = retime_s1_45_reg_reg_IQ;
 reg retime_s1_93_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_93_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_93_reg_reg_IQ <= mul_22_25_n_1454;
     end
 assign n_55 = retime_s1_93_reg_reg_IQ;
 reg retime_s1_46_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_46_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_46_reg_reg_IQ <= mul_22_25_n_1362;
     end
 assign n_107 = retime_s1_46_reg_reg_IQ;
 reg retime_s1_48_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_48_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_48_reg_reg_IQ <= mul_22_25_n_1364;
     end
 assign n_105 = retime_s1_48_reg_reg_IQ;
 reg retime_s1_50_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_50_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_50_reg_reg_IQ <= mul_22_25_n_959;
     end
 assign n_103 = retime_s1_50_reg_reg_IQ;
 reg retime_s1_52_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_52_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_52_reg_reg_IQ <= mul_22_25_n_1548;
     end
 assign n_101 = retime_s1_52_reg_reg_IQ;
 reg retime_s1_56_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_56_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_56_reg_reg_IQ <= mul_22_25_n_1500;
     end
 assign n_97 = retime_s1_56_reg_reg_IQ;
 reg retime_s1_59_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_59_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_59_reg_reg_IQ <= mul_22_25_n_1518;
     end
 assign n_94 = retime_s1_59_reg_reg_IQ;
 reg retime_s1_54_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_54_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_54_reg_reg_IQ <= mul_22_25_n_1532;
     end
 assign n_99 = retime_s1_54_reg_reg_IQ;
 reg retime_s1_58_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_58_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_58_reg_reg_IQ <= mul_22_25_n_1003;
     end
 assign n_95 = retime_s1_58_reg_reg_IQ;
 reg retime_s1_62_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_62_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_62_reg_reg_IQ <= mul_22_25_n_1422;
     end
 assign n_91 = retime_s1_62_reg_reg_IQ;
 reg retime_s1_63_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_63_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_63_reg_reg_IQ <= mul_22_25_n_1389;
     end
 assign n_90 = retime_s1_63_reg_reg_IQ;
 reg retime_s1_65_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_65_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_65_reg_reg_IQ <= mul_22_25_n_1486;
     end
 assign n_88 = retime_s1_65_reg_reg_IQ;
 reg retime_s1_66_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_66_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_66_reg_reg_IQ <= mul_22_25_n_1406;
     end
 assign n_87 = retime_s1_66_reg_reg_IQ;
 reg retime_s1_67_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_67_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_67_reg_reg_IQ <= mul_22_25_n_1502;
     end
 assign n_86 = retime_s1_67_reg_reg_IQ;
 reg retime_s1_21_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_21_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_21_reg_reg_IQ <= mul_22_25_n_1630;
     end
 assign n_132 = retime_s1_21_reg_reg_IQ;
 reg retime_s1_68_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_68_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_68_reg_reg_IQ <= mul_22_25_n_1598;
     end
 assign n_85 = retime_s1_68_reg_reg_IQ;
 reg retime_s1_72_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_72_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_72_reg_reg_IQ <= mul_22_25_n_1420;
     end
 assign n_81 = retime_s1_72_reg_reg_IQ;
 reg retime_s1_73_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_73_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_73_reg_reg_IQ <= mul_22_25_n_1391;
     end
 assign n_80 = retime_s1_73_reg_reg_IQ;
 reg retime_s1_70_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_70_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_70_reg_reg_IQ <= mul_22_25_n_1534;
     end
 assign n_83 = retime_s1_70_reg_reg_IQ;
 reg retime_s1_74_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_74_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_74_reg_reg_IQ <= mul_22_25_n_984;
     end
 assign n_79 = retime_s1_74_reg_reg_IQ;
 reg retime_s1_71_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_71_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_71_reg_reg_IQ <= mul_22_25_n_1404;
     end
 assign n_82 = retime_s1_71_reg_reg_IQ;
 reg retime_s1_85_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_85_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_85_reg_reg_IQ <= mul_22_25_n_1614;
     end
 assign n_64 = retime_s1_85_reg_reg_IQ;
 reg retime_s1_78_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_78_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_78_reg_reg_IQ <= mul_22_25_n_1004;
     end
 assign n_75 = retime_s1_78_reg_reg_IQ;
 reg retime_s1_80_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_80_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_80_reg_reg_IQ <= mul_22_25_n_1438;
     end
 assign n_73 = retime_s1_80_reg_reg_IQ;
 reg retime_s1_83_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_83_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_83_reg_reg_IQ <= mul_22_25_n_961;
     end
 assign n_69 = retime_s1_83_reg_reg_IQ;
 reg retime_s1_84_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_84_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_84_reg_reg_IQ <= mul_22_25_n_1013;
     end
 assign n_68 = retime_s1_84_reg_reg_IQ;
 reg retime_s1_88_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_88_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_88_reg_reg_IQ <= mul_22_25_n_1015;
     end
 assign n_61 = retime_s1_88_reg_reg_IQ;
 reg retime_s1_89_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_89_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_89_reg_reg_IQ <= mul_22_25_n_1436;
     end
 assign n_60 = retime_s1_89_reg_reg_IQ;
 reg retime_s1_91_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_91_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_91_reg_reg_IQ <= mul_22_25_n_1111;
     end
 assign n_58 = retime_s1_91_reg_reg_IQ;
 reg retime_s1_92_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_92_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_92_reg_reg_IQ <= mul_22_25_n_1011;
     end
 assign n_57 = retime_s1_92_reg_reg_IQ;
 reg retime_s1_86_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_86_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_86_reg_reg_IQ <= mul_22_25_n_979;
     end
 assign n_63 = retime_s1_86_reg_reg_IQ;
 reg retime_s1_76_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_76_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_76_reg_reg_IQ <= mul_22_25_n_1008;
     end
 assign n_77 = retime_s1_76_reg_reg_IQ;
 reg retime_s1_99_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_99_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_99_reg_reg_IQ <= mul_22_25_n_9;
     end
 assign n_45 = retime_s1_99_reg_reg_IQ;
 reg retime_s1_69_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_69_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_69_reg_reg_IQ <= mul_22_25_n_1582;
     end
 assign n_84 = retime_s1_69_reg_reg_IQ;
 reg retime_s1_2_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_2_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_2_reg_reg_IQ <= mul_22_25_n_1352;
     end
 assign n_151 = retime_s1_2_reg_reg_IQ;
 reg retime_s1_4_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_4_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_4_reg_reg_IQ <= mul_22_25_n_1350;
     end
 assign n_149 = retime_s1_4_reg_reg_IQ;
 reg retime_s1_8_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_8_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_8_reg_reg_IQ <= mul_22_25_n_955;
     end
 assign n_145 = retime_s1_8_reg_reg_IQ;
 reg retime_s1_10_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_10_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_10_reg_reg_IQ <= mul_22_25_n_1484;
     end
 assign n_143 = retime_s1_10_reg_reg_IQ;
 reg retime_s1_12_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_12_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_12_reg_reg_IQ <= mul_22_25_n_1468;
     end
 assign n_141 = retime_s1_12_reg_reg_IQ;
 reg retime_s1_15_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_15_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_15_reg_reg_IQ <= mul_22_25_n_960;
     end
 assign n_138 = retime_s1_15_reg_reg_IQ;
 reg retime_s1_16_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_16_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_16_reg_reg_IQ <= mul_22_25_n_1452;
     end
 assign n_137 = retime_s1_16_reg_reg_IQ;
 reg retime_s1_19_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_19_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_19_reg_reg_IQ <= mul_22_25_n_1516;
     end
 assign n_134 = retime_s1_19_reg_reg_IQ;
 reg retime_s1_27_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_27_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_27_reg_reg_IQ <= mul_22_25_n_1612;
     end
 assign n_126 = retime_s1_27_reg_reg_IQ;
 reg retime_s1_94_reg_reg_IQ;
 wire retime_s1_94_reg_reg_IQN;
 assign retime_s1_94_reg_reg_IQN = !retime_s1_94_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_94_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_94_reg_reg_IQ <= mul_22_25_n_1758;
     end
 assign mul_22_25_n_1059 = retime_s1_94_reg_reg_IQN;
 assign mul_22_25_n_1283 = ((mul_22_25_n_687 & mul_22_25_n_513) | (mul_22_25_n_529 & (mul_22_25_n_687
    ^ mul_22_25_n_513)));
 assign mul_22_25_n_1282 = (mul_22_25_n_529 ^ (mul_22_25_n_687 ^ mul_22_25_n_513));
 assign mul_22_25_n_1785 = ((mul_22_25_n_798 & mul_22_25_n_672) | (mul_22_25_n_893 & (mul_22_25_n_798
    ^ mul_22_25_n_672)));
 assign mul_22_25_n_1281 = (mul_22_25_n_893 ^ (mul_22_25_n_798 ^ mul_22_25_n_672));
 assign mul_22_25_n_1746 = ((mul_22_25_n_526 & mul_22_25_n_510) | (mul_22_25_n_714 & (mul_22_25_n_526
    ^ mul_22_25_n_510)));
 assign mul_22_25_n_1747 = (mul_22_25_n_714 ^ (mul_22_25_n_526 ^ mul_22_25_n_510));
 assign mul_22_25_n_1280 = ((mul_22_25_n_885 & mul_22_25_n_649) | (mul_22_25_n_1747 & (mul_22_25_n_885
    ^ mul_22_25_n_649)));
 assign mul_22_25_n_1279 = (mul_22_25_n_1747 ^ (mul_22_25_n_885 ^ mul_22_25_n_649));
 assign mul_22_25_n_1744 = ((mul_22_25_n_622 & mul_22_25_n_797) | (mul_22_25_n_658 & (mul_22_25_n_622
    ^ mul_22_25_n_797)));
 assign mul_22_25_n_1745 = (mul_22_25_n_658 ^ (mul_22_25_n_622 ^ mul_22_25_n_797));
 assign mul_22_25_n_1278 = ((mul_22_25_n_1746 & mul_22_25_n_891) | (mul_22_25_n_1745 & (mul_22_25_n_1746
    ^ mul_22_25_n_891)));
 assign mul_22_25_n_1277 = (mul_22_25_n_1745 ^ (mul_22_25_n_1746 ^ mul_22_25_n_891));
 assign mul_22_25_n_1741 = ((mul_22_25_n_525 & mul_22_25_n_508) | (mul_22_25_n_684 & (mul_22_25_n_525
    ^ mul_22_25_n_508)));
 assign mul_22_25_n_1743 = (mul_22_25_n_684 ^ (mul_22_25_n_525 ^ mul_22_25_n_508));
 assign mul_22_25_n_1739 = ((mul_22_25_n_591 & mul_22_25_n_594) | (mul_22_25_n_888 & (mul_22_25_n_591
    ^ mul_22_25_n_594)));
 assign mul_22_25_n_1742 = (mul_22_25_n_888 ^ (mul_22_25_n_591 ^ mul_22_25_n_594));
 assign mul_22_25_n_1786 = ((mul_22_25_n_1743 & mul_22_25_n_1744) | (mul_22_25_n_1742 & (mul_22_25_n_1743
    ^ mul_22_25_n_1744)));
 assign mul_22_25_n_1276 = (mul_22_25_n_1742 ^ (mul_22_25_n_1743 ^ mul_22_25_n_1744));
 assign mul_22_25_n_1737 = ((mul_22_25_n_795 & mul_22_25_n_578) | (mul_22_25_n_527 & (mul_22_25_n_795
    ^ mul_22_25_n_578)));
 assign mul_22_25_n_1740 = (mul_22_25_n_527 ^ (mul_22_25_n_795 ^ mul_22_25_n_578));
 assign mul_22_25_n_1734 = ((mul_22_25_n_896 & mul_22_25_n_562) | (mul_22_25_n_1741 & (mul_22_25_n_896
    ^ mul_22_25_n_562)));
 assign mul_22_25_n_1738 = (mul_22_25_n_1741 ^ (mul_22_25_n_896 ^ mul_22_25_n_562));
 assign mul_22_25_n_1273 = ((mul_22_25_n_1739 & mul_22_25_n_1740) | (mul_22_25_n_1738 & (mul_22_25_n_1739
    ^ mul_22_25_n_1740)));
 assign mul_22_25_n_1748 = (mul_22_25_n_1738 ^ (mul_22_25_n_1739 ^ mul_22_25_n_1740));
 assign mul_22_25_n_1732 = ((mul_22_25_n_777 & mul_22_25_n_511) | (mul_22_25_n_774 & (mul_22_25_n_777
    ^ mul_22_25_n_511)));
 assign mul_22_25_n_1736 = (mul_22_25_n_774 ^ (mul_22_25_n_777 ^ mul_22_25_n_511));
 assign mul_22_25_n_1731 = ((mul_22_25_n_554 & mul_22_25_n_768) | (mul_22_25_n_762 & (mul_22_25_n_554
    ^ mul_22_25_n_768)));
 assign mul_22_25_n_1735 = (mul_22_25_n_762 ^ (mul_22_25_n_554 ^ mul_22_25_n_768));
 assign mul_22_25_n_1727 = ((mul_22_25_n_1737 & mul_22_25_n_884) | (mul_22_25_n_1736 & (mul_22_25_n_1737
    ^ mul_22_25_n_884)));
 assign mul_22_25_n_1733 = (mul_22_25_n_1736 ^ (mul_22_25_n_1737 ^ mul_22_25_n_884));
 assign mul_22_25_n_1272 = ((mul_22_25_n_1734 & mul_22_25_n_1735) | (mul_22_25_n_1733 & (mul_22_25_n_1734
    ^ mul_22_25_n_1735)));
 assign mul_22_25_n_1749 = (mul_22_25_n_1733 ^ (mul_22_25_n_1734 ^ mul_22_25_n_1735));
 assign mul_22_25_n_1726 = ((mul_22_25_n_642 & mul_22_25_n_616) | (mul_22_25_n_528 & (mul_22_25_n_642
    ^ mul_22_25_n_616)));
 assign mul_22_25_n_1730 = (mul_22_25_n_528 ^ (mul_22_25_n_642 ^ mul_22_25_n_616));
 assign mul_22_25_n_1723 = ((mul_22_25_n_728 & mul_22_25_n_800) | (mul_22_25_n_905 & (mul_22_25_n_728
    ^ mul_22_25_n_800)));
 assign mul_22_25_n_1729 = (mul_22_25_n_905 ^ (mul_22_25_n_728 ^ mul_22_25_n_800));
 assign mul_22_25_n_1721 = ((mul_22_25_n_1731 & mul_22_25_n_1732) | (mul_22_25_n_1730 & (mul_22_25_n_1731
    ^ mul_22_25_n_1732)));
 assign mul_22_25_n_1728 = (mul_22_25_n_1730 ^ (mul_22_25_n_1731 ^ mul_22_25_n_1732));
 assign mul_22_25_n_1271 = ((mul_22_25_n_1728 & mul_22_25_n_1729) | (mul_22_25_n_1727 & (mul_22_25_n_1728
    ^ mul_22_25_n_1729)));
 assign mul_22_25_n_1750 = (mul_22_25_n_1727 ^ (mul_22_25_n_1728 ^ mul_22_25_n_1729));
 assign mul_22_25_n_1719 = ((mul_22_25_n_747 & mul_22_25_n_509) | (mul_22_25_n_789 & (mul_22_25_n_747
    ^ mul_22_25_n_509)));
 assign mul_22_25_n_1724 = (mul_22_25_n_789 ^ (mul_22_25_n_747 ^ mul_22_25_n_509));
 assign mul_22_25_n_1718 = ((mul_22_25_n_522 & mul_22_25_n_816) | (mul_22_25_n_820 & (mul_22_25_n_522
    ^ mul_22_25_n_816)));
 assign mul_22_25_n_1725 = (mul_22_25_n_820 ^ (mul_22_25_n_522 ^ mul_22_25_n_816));
 assign mul_22_25_n_1715 = ((mul_22_25_n_881 & mul_22_25_n_724) | (mul_22_25_n_1726 & (mul_22_25_n_881
    ^ mul_22_25_n_724)));
 assign mul_22_25_n_1722 = (mul_22_25_n_1726 ^ (mul_22_25_n_881 ^ mul_22_25_n_724));
 assign mul_22_25_n_1713 = ((mul_22_25_n_1724 & mul_22_25_n_1725) | (mul_22_25_n_1723 & (mul_22_25_n_1724
    ^ mul_22_25_n_1725)));
 assign mul_22_25_n_1720 = (mul_22_25_n_1723 ^ (mul_22_25_n_1724 ^ mul_22_25_n_1725));
 assign mul_22_25_n_1787 = ((mul_22_25_n_1721 & mul_22_25_n_1722) | (mul_22_25_n_1720 & (mul_22_25_n_1721
    ^ mul_22_25_n_1722)));
 assign mul_22_25_n_1751 = (mul_22_25_n_1720 ^ (mul_22_25_n_1721 ^ mul_22_25_n_1722));
 assign mul_22_25_n_1711 = ((mul_22_25_n_662 & mul_22_25_n_698) | (mul_22_25_n_703 & (mul_22_25_n_662
    ^ mul_22_25_n_698)));
 assign mul_22_25_n_1716 = (mul_22_25_n_703 ^ (mul_22_25_n_662 ^ mul_22_25_n_698));
 assign mul_22_25_n_1710 = ((mul_22_25_n_737 & mul_22_25_n_582) | (mul_22_25_n_802 & (mul_22_25_n_737
    ^ mul_22_25_n_582)));
 assign mul_22_25_n_1717 = (mul_22_25_n_802 ^ (mul_22_25_n_737 ^ mul_22_25_n_582));
 assign mul_22_25_n_1706 = ((mul_22_25_n_1719 & mul_22_25_n_895) | (mul_22_25_n_1718 & (mul_22_25_n_1719
    ^ mul_22_25_n_895)));
 assign mul_22_25_n_1714 = (mul_22_25_n_1718 ^ (mul_22_25_n_1719 ^ mul_22_25_n_895));
 assign mul_22_25_n_1703 = ((mul_22_25_n_1716 & mul_22_25_n_1717) | (mul_22_25_n_1715 & (mul_22_25_n_1716
    ^ mul_22_25_n_1717)));
 assign mul_22_25_n_1712 = (mul_22_25_n_1715 ^ (mul_22_25_n_1716 ^ mul_22_25_n_1717));
 assign mul_22_25_n_1788 = ((mul_22_25_n_1713 & mul_22_25_n_1714) | (mul_22_25_n_1712 & (mul_22_25_n_1713
    ^ mul_22_25_n_1714)));
 assign mul_22_25_n_1752 = (mul_22_25_n_1712 ^ (mul_22_25_n_1713 ^ mul_22_25_n_1714));
 assign mul_22_25_n_1702 = ((mul_22_25_n_530 & mul_22_25_n_506) | (mul_22_25_n_761 & (mul_22_25_n_530
    ^ mul_22_25_n_506)));
 assign mul_22_25_n_1709 = (mul_22_25_n_761 ^ (mul_22_25_n_530 ^ mul_22_25_n_506));
 assign mul_22_25_n_1701 = ((mul_22_25_n_613 & mul_22_25_n_682) | (mul_22_25_n_735 & (mul_22_25_n_613
    ^ mul_22_25_n_682)));
 assign mul_22_25_n_1708 = (mul_22_25_n_735 ^ (mul_22_25_n_613 ^ mul_22_25_n_682));
 assign mul_22_25_n_1698 = ((mul_22_25_n_647 & mul_22_25_n_595) | (mul_22_25_n_883 & (mul_22_25_n_647
    ^ mul_22_25_n_595)));
 assign mul_22_25_n_1707 = (mul_22_25_n_883 ^ (mul_22_25_n_647 ^ mul_22_25_n_595));
 assign mul_22_25_n_1696 = ((mul_22_25_n_1710 & mul_22_25_n_1711) | (mul_22_25_n_1709 & (mul_22_25_n_1710
    ^ mul_22_25_n_1711)));
 assign mul_22_25_n_1705 = (mul_22_25_n_1709 ^ (mul_22_25_n_1710 ^ mul_22_25_n_1711));
 assign mul_22_25_n_1694 = ((mul_22_25_n_1707 & mul_22_25_n_1708) | (mul_22_25_n_1706 & (mul_22_25_n_1707
    ^ mul_22_25_n_1708)));
 assign mul_22_25_n_1704 = (mul_22_25_n_1706 ^ (mul_22_25_n_1707 ^ mul_22_25_n_1708));
 assign mul_22_25_n_1789 = ((mul_22_25_n_1704 & mul_22_25_n_1705) | (mul_22_25_n_1703 & (mul_22_25_n_1704
    ^ mul_22_25_n_1705)));
 assign mul_22_25_n_1753 = (mul_22_25_n_1703 ^ (mul_22_25_n_1704 ^ mul_22_25_n_1705));
 assign mul_22_25_n_1692 = ((mul_22_25_n_801 & mul_22_25_n_828) | (mul_22_25_n_727 & (mul_22_25_n_801
    ^ mul_22_25_n_828)));
 assign mul_22_25_n_1699 = (mul_22_25_n_727 ^ (mul_22_25_n_801 ^ mul_22_25_n_828));
 assign mul_22_25_n_1691 = ((mul_22_25_n_579 & mul_22_25_n_718) | (mul_22_25_n_617 & (mul_22_25_n_579
    ^ mul_22_25_n_718)));
 assign mul_22_25_n_1700 = (mul_22_25_n_617 ^ (mul_22_25_n_579 ^ mul_22_25_n_718));
 assign mul_22_25_n_1687 = ((mul_22_25_n_890 & mul_22_25_n_627) | (mul_22_25_n_1702 & (mul_22_25_n_890
    ^ mul_22_25_n_627)));
 assign mul_22_25_n_1697 = (mul_22_25_n_1702 ^ (mul_22_25_n_890 ^ mul_22_25_n_627));
 assign mul_22_25_n_1685 = ((mul_22_25_n_1700 & mul_22_25_n_1701) | (mul_22_25_n_1699 & (mul_22_25_n_1700
    ^ mul_22_25_n_1701)));
 assign mul_22_25_n_1695 = (mul_22_25_n_1699 ^ (mul_22_25_n_1700 ^ mul_22_25_n_1701));
 assign mul_22_25_n_1683 = ((mul_22_25_n_1697 & mul_22_25_n_1698) | (mul_22_25_n_1696 & (mul_22_25_n_1697
    ^ mul_22_25_n_1698)));
 assign mul_22_25_n_1693 = (mul_22_25_n_1696 ^ (mul_22_25_n_1697 ^ mul_22_25_n_1698));
 assign mul_22_25_n_1790 = ((mul_22_25_n_1694 & mul_22_25_n_1695) | (mul_22_25_n_1693 & (mul_22_25_n_1694
    ^ mul_22_25_n_1695)));
 assign mul_22_25_n_1754 = (mul_22_25_n_1693 ^ (mul_22_25_n_1694 ^ mul_22_25_n_1695));
 assign mul_22_25_n_1681 = ((mul_22_25_n_524 & mul_22_25_n_507) | (mul_22_25_n_601 & (mul_22_25_n_524
    ^ mul_22_25_n_507)));
 assign mul_22_25_n_1689 = (mul_22_25_n_601 ^ (mul_22_25_n_524 ^ mul_22_25_n_507));
 assign mul_22_25_n_1679 = ((mul_22_25_n_821 & mul_22_25_n_598) | (mul_22_25_n_597 & (mul_22_25_n_821
    ^ mul_22_25_n_598)));
 assign mul_22_25_n_1688 = (mul_22_25_n_597 ^ (mul_22_25_n_821 ^ mul_22_25_n_598));
 assign mul_22_25_n_1680 = ((mul_22_25_n_565 & mul_22_25_n_593) | (mul_22_25_n_589 & (mul_22_25_n_565
    ^ mul_22_25_n_593)));
 assign mul_22_25_n_1690 = (mul_22_25_n_589 ^ (mul_22_25_n_565 ^ mul_22_25_n_593));
 assign mul_22_25_n_1675 = ((mul_22_25_n_1692 & mul_22_25_n_882) | (mul_22_25_n_1691 & (mul_22_25_n_1692
    ^ mul_22_25_n_882)));
 assign mul_22_25_n_1686 = (mul_22_25_n_1691 ^ (mul_22_25_n_1692 ^ mul_22_25_n_882));
 assign mul_22_25_n_1673 = ((mul_22_25_n_1689 & mul_22_25_n_1690) | (mul_22_25_n_1688 & (mul_22_25_n_1689
    ^ mul_22_25_n_1690)));
 assign mul_22_25_n_1684 = (mul_22_25_n_1688 ^ (mul_22_25_n_1689 ^ mul_22_25_n_1690));
 assign mul_22_25_n_1671 = ((mul_22_25_n_1686 & mul_22_25_n_1687) | (mul_22_25_n_1685 & (mul_22_25_n_1686
    ^ mul_22_25_n_1687)));
 assign mul_22_25_n_1682 = (mul_22_25_n_1685 ^ (mul_22_25_n_1686 ^ mul_22_25_n_1687));
 assign mul_22_25_n_1791 = ((mul_22_25_n_1683 & mul_22_25_n_1684) | (mul_22_25_n_1682 & (mul_22_25_n_1683
    ^ mul_22_25_n_1684)));
 assign mul_22_25_n_1755 = (mul_22_25_n_1682 ^ (mul_22_25_n_1683 ^ mul_22_25_n_1684));
 assign mul_22_25_n_1669 = ((mul_22_25_n_574 & mul_22_25_n_739) | (mul_22_25_n_794 & (mul_22_25_n_574
    ^ mul_22_25_n_739)));
 assign mul_22_25_n_1678 = (mul_22_25_n_794 ^ (mul_22_25_n_574 ^ mul_22_25_n_739));
 assign mul_22_25_n_1668 = ((mul_22_25_n_630 & mul_22_25_n_568) | (mul_22_25_n_644 & (mul_22_25_n_630
    ^ mul_22_25_n_568)));
 assign mul_22_25_n_1677 = (mul_22_25_n_644 ^ (mul_22_25_n_630 ^ mul_22_25_n_568));
 assign mul_22_25_n_1664 = ((mul_22_25_n_577 & mul_22_25_n_564) | (mul_22_25_n_892 & (mul_22_25_n_577
    ^ mul_22_25_n_564)));
 assign mul_22_25_n_1676 = (mul_22_25_n_892 ^ (mul_22_25_n_577 ^ mul_22_25_n_564));
 assign mul_22_25_n_1662 = ((mul_22_25_n_1680 & mul_22_25_n_1681) | (mul_22_25_n_1679 & (mul_22_25_n_1680
    ^ mul_22_25_n_1681)));
 assign mul_22_25_n_1674 = (mul_22_25_n_1679 ^ (mul_22_25_n_1680 ^ mul_22_25_n_1681));
 assign mul_22_25_n_1661 = ((mul_22_25_n_1677 & mul_22_25_n_1678) | (mul_22_25_n_1676 & (mul_22_25_n_1677
    ^ mul_22_25_n_1678)));
 assign mul_22_25_n_1672 = (mul_22_25_n_1676 ^ (mul_22_25_n_1677 ^ mul_22_25_n_1678));
 assign mul_22_25_n_1658 = ((mul_22_25_n_1674 & mul_22_25_n_1675) | (mul_22_25_n_1673 & (mul_22_25_n_1674
    ^ mul_22_25_n_1675)));
 assign mul_22_25_n_1670 = (mul_22_25_n_1673 ^ (mul_22_25_n_1674 ^ mul_22_25_n_1675));
 assign mul_22_25_n_1792 = ((mul_22_25_n_1671 & mul_22_25_n_1672) | (mul_22_25_n_1670 & (mul_22_25_n_1671
    ^ mul_22_25_n_1672)));
 assign mul_22_25_n_1756 = (mul_22_25_n_1670 ^ (mul_22_25_n_1671 ^ mul_22_25_n_1672));
 assign mul_22_25_n_1656 = ((mul_22_25_n_543 & mul_22_25_n_512) | (mul_22_25_n_775 & (mul_22_25_n_543
    ^ mul_22_25_n_512)));
 assign mul_22_25_n_1666 = (mul_22_25_n_775 ^ (mul_22_25_n_543 ^ mul_22_25_n_512));
 assign mul_22_25_n_1655 = ((mul_22_25_n_769 & mul_22_25_n_822) | (mul_22_25_n_722 & (mul_22_25_n_769
    ^ mul_22_25_n_822)));
 assign mul_22_25_n_1665 = (mul_22_25_n_722 ^ (mul_22_25_n_769 ^ mul_22_25_n_822));
 assign mul_22_25_n_1654 = ((mul_22_25_n_765 & mul_22_25_n_756) | (mul_22_25_n_784 & (mul_22_25_n_765
    ^ mul_22_25_n_756)));
 assign mul_22_25_n_1667 = (mul_22_25_n_784 ^ (mul_22_25_n_765 ^ mul_22_25_n_756));
 assign mul_22_25_n_1650 = ((mul_22_25_n_887 & mul_22_25_n_760) | (mul_22_25_n_1669 & (mul_22_25_n_887
    ^ mul_22_25_n_760)));
 assign mul_22_25_n_1663 = (mul_22_25_n_1669 ^ (mul_22_25_n_887 ^ mul_22_25_n_760));
 assign mul_22_25_n_1648 = ((mul_22_25_n_1667 & mul_22_25_n_1668) | (mul_22_25_n_1666 & (mul_22_25_n_1667
    ^ mul_22_25_n_1668)));
 assign mul_22_25_n_1660 = (mul_22_25_n_1666 ^ (mul_22_25_n_1667 ^ mul_22_25_n_1668));
 assign mul_22_25_n_1646 = ((mul_22_25_n_1664 & mul_22_25_n_1665) | (mul_22_25_n_1663 & (mul_22_25_n_1664
    ^ mul_22_25_n_1665)));
 assign mul_22_25_n_1659 = (mul_22_25_n_1663 ^ (mul_22_25_n_1664 ^ mul_22_25_n_1665));
 assign mul_22_25_n_1644 = ((mul_22_25_n_1661 & mul_22_25_n_1662) | (mul_22_25_n_1660 & (mul_22_25_n_1661
    ^ mul_22_25_n_1662)));
 assign mul_22_25_n_1657 = (mul_22_25_n_1660 ^ (mul_22_25_n_1661 ^ mul_22_25_n_1662));
 assign mul_22_25_n_1793 = ((mul_22_25_n_1658 & mul_22_25_n_1659) | (mul_22_25_n_1657 & (mul_22_25_n_1658
    ^ mul_22_25_n_1659)));
 assign mul_22_25_n_1757 = (mul_22_25_n_1657 ^ (mul_22_25_n_1658 ^ mul_22_25_n_1659));
 assign mul_22_25_n_1642 = ((mul_22_25_n_638 & mul_22_25_n_689) | (mul_22_25_n_643 & (mul_22_25_n_638
    ^ mul_22_25_n_689)));
 assign mul_22_25_n_1652 = (mul_22_25_n_643 ^ (mul_22_25_n_638 ^ mul_22_25_n_689));
 assign mul_22_25_n_1640 = ((mul_22_25_n_799 & mul_22_25_n_688) | (mul_22_25_n_733 & (mul_22_25_n_799
    ^ mul_22_25_n_688)));
 assign mul_22_25_n_1651 = (mul_22_25_n_733 ^ (mul_22_25_n_799 ^ mul_22_25_n_688));
 assign mul_22_25_n_1641 = ((mul_22_25_n_730 & mul_22_25_n_655) | (mul_22_25_n_583 & (mul_22_25_n_730
    ^ mul_22_25_n_655)));
 assign mul_22_25_n_1653 = (mul_22_25_n_583 ^ (mul_22_25_n_730 ^ mul_22_25_n_655));
 assign mul_22_25_n_1635 = ((mul_22_25_n_1656 & mul_22_25_n_899) | (mul_22_25_n_1655 & (mul_22_25_n_1656
    ^ mul_22_25_n_899)));
 assign mul_22_25_n_1649 = (mul_22_25_n_1655 ^ (mul_22_25_n_1656 ^ mul_22_25_n_899));
 assign mul_22_25_n_1634 = ((mul_22_25_n_1653 & mul_22_25_n_1654) | (mul_22_25_n_1652 & (mul_22_25_n_1653
    ^ mul_22_25_n_1654)));
 assign mul_22_25_n_1647 = (mul_22_25_n_1652 ^ (mul_22_25_n_1653 ^ mul_22_25_n_1654));
 assign mul_22_25_n_1630 = ((mul_22_25_n_1650 & mul_22_25_n_1651) | (mul_22_25_n_1649 & (mul_22_25_n_1650
    ^ mul_22_25_n_1651)));
 assign mul_22_25_n_1645 = (mul_22_25_n_1649 ^ (mul_22_25_n_1650 ^ mul_22_25_n_1651));
 assign mul_22_25_n_1629 = ((mul_22_25_n_1647 & mul_22_25_n_1648) | (mul_22_25_n_1646 & (mul_22_25_n_1647
    ^ mul_22_25_n_1648)));
 assign mul_22_25_n_1643 = (mul_22_25_n_1646 ^ (mul_22_25_n_1647 ^ mul_22_25_n_1648));
 assign mul_22_25_n_1794 = ((mul_22_25_n_1644 & mul_22_25_n_1645) | (mul_22_25_n_1643 & (mul_22_25_n_1644
    ^ mul_22_25_n_1645)));
 assign mul_22_25_n_1758 = (mul_22_25_n_1643 ^ (mul_22_25_n_1644 ^ mul_22_25_n_1645));
 assign mul_22_25_n_1626 = ((mul_22_25_n_544 & mul_22_25_n_514) | (mul_22_25_n_576 & (mul_22_25_n_544
    ^ mul_22_25_n_514)));
 assign mul_22_25_n_1639 = (mul_22_25_n_576 ^ (mul_22_25_n_544 ^ mul_22_25_n_514));
 assign mul_22_25_n_1627 = ((mul_22_25_n_750 & mul_22_25_n_742) | (mul_22_25_n_779 & (mul_22_25_n_750
    ^ mul_22_25_n_742)));
 assign mul_22_25_n_1638 = (mul_22_25_n_779 ^ (mul_22_25_n_750 ^ mul_22_25_n_742));
 assign mul_22_25_n_1625 = ((mul_22_25_n_804 & mul_22_25_n_796) | (mul_22_25_n_621 & (mul_22_25_n_804
    ^ mul_22_25_n_796)));
 assign mul_22_25_n_1637 = (mul_22_25_n_621 ^ (mul_22_25_n_804 ^ mul_22_25_n_796));
 assign mul_22_25_n_1621 = ((mul_22_25_n_819 & mul_22_25_n_817) | (mul_22_25_n_886 & (mul_22_25_n_819
    ^ mul_22_25_n_817)));
 assign mul_22_25_n_1636 = (mul_22_25_n_886 ^ (mul_22_25_n_819 ^ mul_22_25_n_817));
 assign mul_22_25_n_1620 = ((mul_22_25_n_1641 & mul_22_25_n_1642) | (mul_22_25_n_1640 & (mul_22_25_n_1641
    ^ mul_22_25_n_1642)));
 assign mul_22_25_n_1633 = (mul_22_25_n_1640 ^ (mul_22_25_n_1641 ^ mul_22_25_n_1642));
 assign mul_22_25_n_1617 = ((mul_22_25_n_1638 & mul_22_25_n_1639) | (mul_22_25_n_1637 & (mul_22_25_n_1638
    ^ mul_22_25_n_1639)));
 assign mul_22_25_n_1632 = (mul_22_25_n_1637 ^ (mul_22_25_n_1638 ^ mul_22_25_n_1639));
 assign mul_22_25_n_1614 = ((mul_22_25_n_1635 & mul_22_25_n_1636) | (mul_22_25_n_1634 & (mul_22_25_n_1635
    ^ mul_22_25_n_1636)));
 assign mul_22_25_n_1631 = (mul_22_25_n_1634 ^ (mul_22_25_n_1635 ^ mul_22_25_n_1636));
 assign mul_22_25_n_1612 = ((mul_22_25_n_1632 & mul_22_25_n_1633) | (mul_22_25_n_1631 & (mul_22_25_n_1632
    ^ mul_22_25_n_1633)));
 assign mul_22_25_n_1628 = (mul_22_25_n_1631 ^ (mul_22_25_n_1632 ^ mul_22_25_n_1633));
 assign mul_22_25_n_1795 = ((n_113 & n_132) | (n_125 & (n_113 ^ n_132)));
 assign mul_22_25_n_1759 = (n_125 ^ (n_113 ^ n_132));
 assign mul_22_25_n_1610 = ((mul_22_25_n_666 & mul_22_25_n_596) | (mul_22_25_n_700 & (mul_22_25_n_666
    ^ mul_22_25_n_596)));
 assign mul_22_25_n_1623 = (mul_22_25_n_700 ^ (mul_22_25_n_666 ^ mul_22_25_n_596));
 assign mul_22_25_n_1609 = ((mul_22_25_n_585 & mul_22_25_n_743) | (mul_22_25_n_461 & (mul_22_25_n_585
    ^ mul_22_25_n_743)));
 assign mul_22_25_n_1622 = (mul_22_25_n_461 ^ (mul_22_25_n_585 ^ mul_22_25_n_743));
 assign mul_22_25_n_1611 = ((mul_22_25_n_696 & mul_22_25_n_523) | (mul_22_25_n_694 & (mul_22_25_n_696
    ^ mul_22_25_n_523)));
 assign mul_22_25_n_1624 = (mul_22_25_n_694 ^ (mul_22_25_n_696 ^ mul_22_25_n_523));
 assign mul_22_25_n_1605 = ((mul_22_25_n_904 & mul_22_25_n_691) | (mul_22_25_n_1627 & (mul_22_25_n_904
    ^ mul_22_25_n_691)));
 assign mul_22_25_n_1619 = (mul_22_25_n_1627 ^ (mul_22_25_n_904 ^ mul_22_25_n_691));
 assign mul_22_25_n_1603 = ((mul_22_25_n_1625 & mul_22_25_n_1626) | (mul_22_25_n_1624 & (mul_22_25_n_1625
    ^ mul_22_25_n_1626)));
 assign mul_22_25_n_1618 = (mul_22_25_n_1624 ^ (mul_22_25_n_1625 ^ mul_22_25_n_1626));
 assign mul_22_25_n_1601 = ((mul_22_25_n_1622 & mul_22_25_n_1623) | (mul_22_25_n_1621 & (mul_22_25_n_1622
    ^ mul_22_25_n_1623)));
 assign mul_22_25_n_1616 = (mul_22_25_n_1621 ^ (mul_22_25_n_1622 ^ mul_22_25_n_1623));
 assign mul_22_25_n_1599 = ((mul_22_25_n_1619 & mul_22_25_n_1620) | (mul_22_25_n_1618 & (mul_22_25_n_1619
    ^ mul_22_25_n_1620)));
 assign mul_22_25_n_1615 = (mul_22_25_n_1618 ^ (mul_22_25_n_1619 ^ mul_22_25_n_1620));
 assign mul_22_25_n_1596 = ((mul_22_25_n_1616 & mul_22_25_n_1617) | (mul_22_25_n_1615 & (mul_22_25_n_1616
    ^ mul_22_25_n_1617)));
 assign mul_22_25_n_1613 = (mul_22_25_n_1615 ^ (mul_22_25_n_1616 ^ mul_22_25_n_1617));
 assign mul_22_25_n_1796 = ((n_123 & n_64) | (n_126 & (n_123 ^ n_64)));
 assign mul_22_25_n_1760 = (n_126 ^ (n_123 ^ n_64));
 assign mul_22_25_n_1594 = ((mul_22_25_n_675 & mul_22_25_n_678) | (mul_22_25_n_674 & (mul_22_25_n_675
    ^ mul_22_25_n_678)));
 assign mul_22_25_n_1608 = (mul_22_25_n_674 ^ (mul_22_25_n_675 ^ mul_22_25_n_678));
 assign mul_22_25_n_1593 = ((mul_22_25_n_667 & mul_22_25_n_776) | (mul_22_25_n_473 & (mul_22_25_n_667
    ^ mul_22_25_n_776)));
 assign mul_22_25_n_1607 = (mul_22_25_n_473 ^ (mul_22_25_n_667 ^ mul_22_25_n_776));
 assign mul_22_25_n_1595 = ((mul_22_25_n_633 & mul_22_25_n_771) | (mul_22_25_n_757 & (mul_22_25_n_633
    ^ mul_22_25_n_771)));
 assign mul_22_25_n_1606 = (mul_22_25_n_757 ^ (mul_22_25_n_633 ^ mul_22_25_n_771));
 assign mul_22_25_n_1589 = ((mul_22_25_n_880 & mul_22_25_n_903) | (mul_22_25_n_1611 & (mul_22_25_n_880
    ^ mul_22_25_n_903)));
 assign mul_22_25_n_1604 = (mul_22_25_n_1611 ^ (mul_22_25_n_880 ^ mul_22_25_n_903));
 assign mul_22_25_n_1587 = ((mul_22_25_n_1609 & mul_22_25_n_1610) | (mul_22_25_n_1608 & (mul_22_25_n_1609
    ^ mul_22_25_n_1610)));
 assign mul_22_25_n_1602 = (mul_22_25_n_1608 ^ (mul_22_25_n_1609 ^ mul_22_25_n_1610));
 assign mul_22_25_n_1584 = ((mul_22_25_n_1606 & mul_22_25_n_1607) | (mul_22_25_n_1605 & (mul_22_25_n_1606
    ^ mul_22_25_n_1607)));
 assign mul_22_25_n_1600 = (mul_22_25_n_1605 ^ (mul_22_25_n_1606 ^ mul_22_25_n_1607));
 assign mul_22_25_n_1583 = ((mul_22_25_n_1603 & mul_22_25_n_1604) | (mul_22_25_n_1602 & (mul_22_25_n_1603
    ^ mul_22_25_n_1604)));
 assign mul_22_25_n_1598 = (mul_22_25_n_1602 ^ (mul_22_25_n_1603 ^ mul_22_25_n_1604));
 assign mul_22_25_n_1580 = ((mul_22_25_n_1600 & mul_22_25_n_1601) | (mul_22_25_n_1599 & (mul_22_25_n_1600
    ^ mul_22_25_n_1601)));
 assign mul_22_25_n_1597 = (mul_22_25_n_1599 ^ (mul_22_25_n_1600 ^ mul_22_25_n_1601));
 assign mul_22_25_n_1797 = ((n_121 & n_85) | (n_124 & (n_121 ^ n_85)));
 assign mul_22_25_n_1761 = (n_124 ^ (n_121 ^ n_85));
 assign mul_22_25_n_1578 = ((mul_22_25_n_653 & mul_22_25_n_720) | (mul_22_25_n_690 & (mul_22_25_n_653
    ^ mul_22_25_n_720)));
 assign mul_22_25_n_1592 = (mul_22_25_n_690 ^ (mul_22_25_n_653 ^ mul_22_25_n_720));
 assign mul_22_25_n_1577 = ((mul_22_25_n_600 & mul_22_25_n_612) | (mul_22_25_n_495 & (mul_22_25_n_600
    ^ mul_22_25_n_612)));
 assign mul_22_25_n_1591 = (mul_22_25_n_495 ^ (mul_22_25_n_600 ^ mul_22_25_n_612));
 assign mul_22_25_n_1579 = ((mul_22_25_n_715 & mul_22_25_n_826) | (mul_22_25_n_778 & (mul_22_25_n_715
    ^ mul_22_25_n_826)));
 assign mul_22_25_n_1590 = (mul_22_25_n_778 ^ (mul_22_25_n_715 ^ mul_22_25_n_826));
 assign mul_22_25_n_1573 = ((mul_22_25_n_877 & mul_22_25_n_902) | (mul_22_25_n_1595 & (mul_22_25_n_877
    ^ mul_22_25_n_902)));
 assign mul_22_25_n_1588 = (mul_22_25_n_1595 ^ (mul_22_25_n_877 ^ mul_22_25_n_902));
 assign mul_22_25_n_1571 = ((mul_22_25_n_1593 & mul_22_25_n_1594) | (mul_22_25_n_1592 & (mul_22_25_n_1593
    ^ mul_22_25_n_1594)));
 assign mul_22_25_n_1586 = (mul_22_25_n_1592 ^ (mul_22_25_n_1593 ^ mul_22_25_n_1594));
 assign mul_22_25_n_1568 = ((mul_22_25_n_1590 & mul_22_25_n_1591) | (mul_22_25_n_1589 & (mul_22_25_n_1590
    ^ mul_22_25_n_1591)));
 assign mul_22_25_n_1585 = (mul_22_25_n_1589 ^ (mul_22_25_n_1590 ^ mul_22_25_n_1591));
 assign mul_22_25_n_1567 = ((mul_22_25_n_1587 & mul_22_25_n_1588) | (mul_22_25_n_1586 & (mul_22_25_n_1587
    ^ mul_22_25_n_1588)));
 assign mul_22_25_n_1582 = (mul_22_25_n_1586 ^ (mul_22_25_n_1587 ^ mul_22_25_n_1588));
 assign mul_22_25_n_1564 = ((mul_22_25_n_1584 & mul_22_25_n_1585) | (mul_22_25_n_1583 & (mul_22_25_n_1584
    ^ mul_22_25_n_1585)));
 assign mul_22_25_n_1581 = (mul_22_25_n_1583 ^ (mul_22_25_n_1584 ^ mul_22_25_n_1585));
 assign mul_22_25_n_1798 = ((n_111 & n_84) | (n_122 & (n_111 ^ n_84)));
 assign mul_22_25_n_1762 = (n_122 ^ (n_111 ^ n_84));
 assign mul_22_25_n_1562 = ((mul_22_25_n_751 & mul_22_25_n_602) | (mul_22_25_n_628 & (mul_22_25_n_751
    ^ mul_22_25_n_602)));
 assign mul_22_25_n_1576 = (mul_22_25_n_628 ^ (mul_22_25_n_751 ^ mul_22_25_n_602));
 assign mul_22_25_n_1561 = ((mul_22_25_n_625 & mul_22_25_n_646) | (mul_22_25_n_501 & (mul_22_25_n_625
    ^ mul_22_25_n_646)));
 assign mul_22_25_n_1575 = (mul_22_25_n_501 ^ (mul_22_25_n_625 ^ mul_22_25_n_646));
 assign mul_22_25_n_1563 = ((mul_22_25_n_584 & mul_22_25_n_661) | (mul_22_25_n_620 & (mul_22_25_n_584
    ^ mul_22_25_n_661)));
 assign mul_22_25_n_1574 = (mul_22_25_n_620 ^ (mul_22_25_n_584 ^ mul_22_25_n_661));
 assign mul_22_25_n_1557 = ((mul_22_25_n_870 & mul_22_25_n_901) | (mul_22_25_n_1579 & (mul_22_25_n_870
    ^ mul_22_25_n_901)));
 assign mul_22_25_n_1572 = (mul_22_25_n_1579 ^ (mul_22_25_n_870 ^ mul_22_25_n_901));
 assign mul_22_25_n_1555 = ((mul_22_25_n_1577 & mul_22_25_n_1578) | (mul_22_25_n_1576 & (mul_22_25_n_1577
    ^ mul_22_25_n_1578)));
 assign mul_22_25_n_1570 = (mul_22_25_n_1576 ^ (mul_22_25_n_1577 ^ mul_22_25_n_1578));
 assign mul_22_25_n_1552 = ((mul_22_25_n_1574 & mul_22_25_n_1575) | (mul_22_25_n_1573 & (mul_22_25_n_1574
    ^ mul_22_25_n_1575)));
 assign mul_22_25_n_1569 = (mul_22_25_n_1573 ^ (mul_22_25_n_1574 ^ mul_22_25_n_1575));
 assign mul_22_25_n_1551 = ((mul_22_25_n_1571 & mul_22_25_n_1572) | (mul_22_25_n_1570 & (mul_22_25_n_1571
    ^ mul_22_25_n_1572)));
 assign mul_22_25_n_1566 = (mul_22_25_n_1570 ^ (mul_22_25_n_1571 ^ mul_22_25_n_1572));
 assign mul_22_25_n_1548 = ((mul_22_25_n_1568 & mul_22_25_n_1569) | (mul_22_25_n_1567 & (mul_22_25_n_1568
    ^ mul_22_25_n_1569)));
 assign mul_22_25_n_1565 = (mul_22_25_n_1567 ^ (mul_22_25_n_1568 ^ mul_22_25_n_1569));
 assign mul_22_25_n_1799 = ((n_100 & n_48) | (n_112 & (n_100 ^ n_48)));
 assign mul_22_25_n_1763 = (n_112 ^ (n_100 ^ n_48));
 assign mul_22_25_n_1546 = ((mul_22_25_n_610 & mul_22_25_n_611) | (mul_22_25_n_609 & (mul_22_25_n_610
    ^ mul_22_25_n_611)));
 assign mul_22_25_n_1560 = (mul_22_25_n_609 ^ (mul_22_25_n_610 ^ mul_22_25_n_611));
 assign mul_22_25_n_1545 = ((mul_22_25_n_607 & mul_22_25_n_608) | (mul_22_25_n_477 & (mul_22_25_n_607
    ^ mul_22_25_n_608)));
 assign mul_22_25_n_1559 = (mul_22_25_n_477 ^ (mul_22_25_n_607 ^ mul_22_25_n_608));
 assign mul_22_25_n_1547 = ((mul_22_25_n_605 & mul_22_25_n_780) | (mul_22_25_n_603 & (mul_22_25_n_605
    ^ mul_22_25_n_780)));
 assign mul_22_25_n_1558 = (mul_22_25_n_603 ^ (mul_22_25_n_605 ^ mul_22_25_n_780));
 assign mul_22_25_n_1541 = ((mul_22_25_n_869 & mul_22_25_n_894) | (mul_22_25_n_1563 & (mul_22_25_n_869
    ^ mul_22_25_n_894)));
 assign mul_22_25_n_1556 = (mul_22_25_n_1563 ^ (mul_22_25_n_869 ^ mul_22_25_n_894));
 assign mul_22_25_n_1539 = ((mul_22_25_n_1561 & mul_22_25_n_1562) | (mul_22_25_n_1560 & (mul_22_25_n_1561
    ^ mul_22_25_n_1562)));
 assign mul_22_25_n_1554 = (mul_22_25_n_1560 ^ (mul_22_25_n_1561 ^ mul_22_25_n_1562));
 assign mul_22_25_n_1536 = ((mul_22_25_n_1558 & mul_22_25_n_1559) | (mul_22_25_n_1557 & (mul_22_25_n_1558
    ^ mul_22_25_n_1559)));
 assign mul_22_25_n_1553 = (mul_22_25_n_1557 ^ (mul_22_25_n_1558 ^ mul_22_25_n_1559));
 assign mul_22_25_n_1535 = ((mul_22_25_n_1555 & mul_22_25_n_1556) | (mul_22_25_n_1554 & (mul_22_25_n_1555
    ^ mul_22_25_n_1556)));
 assign mul_22_25_n_1550 = (mul_22_25_n_1554 ^ (mul_22_25_n_1555 ^ mul_22_25_n_1556));
 assign mul_22_25_n_1532 = ((mul_22_25_n_1552 & mul_22_25_n_1553) | (mul_22_25_n_1551 & (mul_22_25_n_1552
    ^ mul_22_25_n_1553)));
 assign mul_22_25_n_1549 = (mul_22_25_n_1551 ^ (mul_22_25_n_1552 ^ mul_22_25_n_1553));
 assign mul_22_25_n_1800 = ((n_98 & n_135) | (n_101 & (n_98 ^ n_135)));
 assign mul_22_25_n_1764 = (n_101 ^ (n_98 ^ n_135));
 assign mul_22_25_n_1530 = ((mul_22_25_n_793 & mul_22_25_n_656) | (mul_22_25_n_592 & (mul_22_25_n_793
    ^ mul_22_25_n_656)));
 assign mul_22_25_n_1544 = (mul_22_25_n_592 ^ (mul_22_25_n_793 ^ mul_22_25_n_656));
 assign mul_22_25_n_1529 = ((mul_22_25_n_588 & mul_22_25_n_590) | (mul_22_25_n_504 & (mul_22_25_n_588
    ^ mul_22_25_n_590)));
 assign mul_22_25_n_1543 = (mul_22_25_n_504 ^ (mul_22_25_n_588 ^ mul_22_25_n_590));
 assign mul_22_25_n_1531 = ((mul_22_25_n_686 & mul_22_25_n_626) | (mul_22_25_n_587 & (mul_22_25_n_686
    ^ mul_22_25_n_626)));
 assign mul_22_25_n_1542 = (mul_22_25_n_587 ^ (mul_22_25_n_686 ^ mul_22_25_n_626));
 assign mul_22_25_n_1525 = ((mul_22_25_n_872 & mul_22_25_n_898) | (mul_22_25_n_1547 & (mul_22_25_n_872
    ^ mul_22_25_n_898)));
 assign mul_22_25_n_1540 = (mul_22_25_n_1547 ^ (mul_22_25_n_872 ^ mul_22_25_n_898));
 assign mul_22_25_n_1523 = ((mul_22_25_n_1545 & mul_22_25_n_1546) | (mul_22_25_n_1544 & (mul_22_25_n_1545
    ^ mul_22_25_n_1546)));
 assign mul_22_25_n_1538 = (mul_22_25_n_1544 ^ (mul_22_25_n_1545 ^ mul_22_25_n_1546));
 assign mul_22_25_n_1520 = ((mul_22_25_n_1542 & mul_22_25_n_1543) | (mul_22_25_n_1541 & (mul_22_25_n_1542
    ^ mul_22_25_n_1543)));
 assign mul_22_25_n_1537 = (mul_22_25_n_1541 ^ (mul_22_25_n_1542 ^ mul_22_25_n_1543));
 assign mul_22_25_n_1519 = ((mul_22_25_n_1539 & mul_22_25_n_1540) | (mul_22_25_n_1538 & (mul_22_25_n_1539
    ^ mul_22_25_n_1540)));
 assign mul_22_25_n_1534 = (mul_22_25_n_1538 ^ (mul_22_25_n_1539 ^ mul_22_25_n_1540));
 assign mul_22_25_n_1516 = ((mul_22_25_n_1536 & mul_22_25_n_1537) | (mul_22_25_n_1535 & (mul_22_25_n_1536
    ^ mul_22_25_n_1537)));
 assign mul_22_25_n_1533 = (mul_22_25_n_1535 ^ (mul_22_25_n_1536 ^ mul_22_25_n_1537));
 assign mul_22_25_n_1801 = ((n_133 & n_83) | (n_99 & (n_133 ^ n_83)));
 assign mul_22_25_n_1765 = (n_99 ^ (n_133 ^ n_83));
 assign mul_22_25_n_1514 = ((mul_22_25_n_573 & mul_22_25_n_575) | (mul_22_25_n_572 & (mul_22_25_n_573
    ^ mul_22_25_n_575)));
 assign mul_22_25_n_1528 = (mul_22_25_n_572 ^ (mul_22_25_n_573 ^ mul_22_25_n_575));
 assign mul_22_25_n_1513 = ((mul_22_25_n_570 & mul_22_25_n_571) | (mul_22_25_n_460 & (mul_22_25_n_570
    ^ mul_22_25_n_571)));
 assign mul_22_25_n_1527 = (mul_22_25_n_460 ^ (mul_22_25_n_570 ^ mul_22_25_n_571));
 assign mul_22_25_n_1515 = ((mul_22_25_n_567 & mul_22_25_n_606) | (mul_22_25_n_566 & (mul_22_25_n_567
    ^ mul_22_25_n_606)));
 assign mul_22_25_n_1526 = (mul_22_25_n_566 ^ (mul_22_25_n_567 ^ mul_22_25_n_606));
 assign mul_22_25_n_1509 = ((mul_22_25_n_873 & mul_22_25_n_897) | (mul_22_25_n_1531 & (mul_22_25_n_873
    ^ mul_22_25_n_897)));
 assign mul_22_25_n_1524 = (mul_22_25_n_1531 ^ (mul_22_25_n_873 ^ mul_22_25_n_897));
 assign mul_22_25_n_1507 = ((mul_22_25_n_1529 & mul_22_25_n_1530) | (mul_22_25_n_1528 & (mul_22_25_n_1529
    ^ mul_22_25_n_1530)));
 assign mul_22_25_n_1522 = (mul_22_25_n_1528 ^ (mul_22_25_n_1529 ^ mul_22_25_n_1530));
 assign mul_22_25_n_1504 = ((mul_22_25_n_1526 & mul_22_25_n_1527) | (mul_22_25_n_1525 & (mul_22_25_n_1526
    ^ mul_22_25_n_1527)));
 assign mul_22_25_n_1521 = (mul_22_25_n_1525 ^ (mul_22_25_n_1526 ^ mul_22_25_n_1527));
 assign mul_22_25_n_1503 = ((mul_22_25_n_1523 & mul_22_25_n_1524) | (mul_22_25_n_1522 & (mul_22_25_n_1523
    ^ mul_22_25_n_1524)));
 assign mul_22_25_n_1518 = (mul_22_25_n_1522 ^ (mul_22_25_n_1523 ^ mul_22_25_n_1524));
 assign mul_22_25_n_1500 = ((mul_22_25_n_1520 & mul_22_25_n_1521) | (mul_22_25_n_1519 & (mul_22_25_n_1520
    ^ mul_22_25_n_1521)));
 assign mul_22_25_n_1517 = (mul_22_25_n_1519 ^ (mul_22_25_n_1520 ^ mul_22_25_n_1521));
 assign mul_22_25_n_1802 = ((n_96 & n_94) | (n_134 & (n_96 ^ n_94)));
 assign mul_22_25_n_1766 = (n_134 ^ (n_96 ^ n_94));
 assign mul_22_25_n_1498 = ((mul_22_25_n_772 & mul_22_25_n_654) | (mul_22_25_n_792 & (mul_22_25_n_772
    ^ mul_22_25_n_654)));
 assign mul_22_25_n_1512 = (mul_22_25_n_792 ^ (mul_22_25_n_772 ^ mul_22_25_n_654));
 assign mul_22_25_n_1497 = ((mul_22_25_n_785 & mul_22_25_n_790) | (mul_22_25_n_476 & (mul_22_25_n_785
    ^ mul_22_25_n_790)));
 assign mul_22_25_n_1511 = (mul_22_25_n_476 ^ (mul_22_25_n_785 ^ mul_22_25_n_790));
 assign mul_22_25_n_1499 = ((mul_22_25_n_782 & mul_22_25_n_783) | (mul_22_25_n_781 & (mul_22_25_n_782
    ^ mul_22_25_n_783)));
 assign mul_22_25_n_1510 = (mul_22_25_n_781 ^ (mul_22_25_n_782 ^ mul_22_25_n_783));
 assign mul_22_25_n_1493 = ((mul_22_25_n_871 & mul_22_25_n_909) | (mul_22_25_n_1515 & (mul_22_25_n_871
    ^ mul_22_25_n_909)));
 assign mul_22_25_n_1508 = (mul_22_25_n_1515 ^ (mul_22_25_n_871 ^ mul_22_25_n_909));
 assign mul_22_25_n_1491 = ((mul_22_25_n_1513 & mul_22_25_n_1514) | (mul_22_25_n_1512 & (mul_22_25_n_1513
    ^ mul_22_25_n_1514)));
 assign mul_22_25_n_1506 = (mul_22_25_n_1512 ^ (mul_22_25_n_1513 ^ mul_22_25_n_1514));
 assign mul_22_25_n_1488 = ((mul_22_25_n_1510 & mul_22_25_n_1511) | (mul_22_25_n_1509 & (mul_22_25_n_1510
    ^ mul_22_25_n_1511)));
 assign mul_22_25_n_1505 = (mul_22_25_n_1509 ^ (mul_22_25_n_1510 ^ mul_22_25_n_1511));
 assign mul_22_25_n_1487 = ((mul_22_25_n_1507 & mul_22_25_n_1508) | (mul_22_25_n_1506 & (mul_22_25_n_1507
    ^ mul_22_25_n_1508)));
 assign mul_22_25_n_1502 = (mul_22_25_n_1506 ^ (mul_22_25_n_1507 ^ mul_22_25_n_1508));
 assign mul_22_25_n_1484 = ((mul_22_25_n_1504 & mul_22_25_n_1505) | (mul_22_25_n_1503 & (mul_22_25_n_1504
    ^ mul_22_25_n_1505)));
 assign mul_22_25_n_1501 = (mul_22_25_n_1503 ^ (mul_22_25_n_1504 ^ mul_22_25_n_1505));
 assign mul_22_25_n_1803 = ((n_142 & n_86) | (n_97 & (n_142 ^ n_86)));
 assign mul_22_25_n_1767 = (n_97 ^ (n_142 ^ n_86));
 assign mul_22_25_n_1482 = ((mul_22_25_n_726 & mul_22_25_n_770) | (mul_22_25_n_719 & (mul_22_25_n_726
    ^ mul_22_25_n_770)));
 assign mul_22_25_n_1496 = (mul_22_25_n_719 ^ (mul_22_25_n_726 ^ mul_22_25_n_770));
 assign mul_22_25_n_1481 = ((mul_22_25_n_740 & mul_22_25_n_734) | (mul_22_25_n_503 & (mul_22_25_n_740
    ^ mul_22_25_n_734)));
 assign mul_22_25_n_1495 = (mul_22_25_n_503 ^ (mul_22_25_n_740 ^ mul_22_25_n_734));
 assign mul_22_25_n_1483 = ((mul_22_25_n_766 & mul_22_25_n_759) | (mul_22_25_n_764 & (mul_22_25_n_766
    ^ mul_22_25_n_759)));
 assign mul_22_25_n_1494 = (mul_22_25_n_764 ^ (mul_22_25_n_766 ^ mul_22_25_n_759));
 assign mul_22_25_n_1477 = ((mul_22_25_n_876 & mul_22_25_n_908) | (mul_22_25_n_1499 & (mul_22_25_n_876
    ^ mul_22_25_n_908)));
 assign mul_22_25_n_1492 = (mul_22_25_n_1499 ^ (mul_22_25_n_876 ^ mul_22_25_n_908));
 assign mul_22_25_n_1475 = ((mul_22_25_n_1497 & mul_22_25_n_1498) | (mul_22_25_n_1496 & (mul_22_25_n_1497
    ^ mul_22_25_n_1498)));
 assign mul_22_25_n_1490 = (mul_22_25_n_1496 ^ (mul_22_25_n_1497 ^ mul_22_25_n_1498));
 assign mul_22_25_n_1472 = ((mul_22_25_n_1494 & mul_22_25_n_1495) | (mul_22_25_n_1493 & (mul_22_25_n_1494
    ^ mul_22_25_n_1495)));
 assign mul_22_25_n_1489 = (mul_22_25_n_1493 ^ (mul_22_25_n_1494 ^ mul_22_25_n_1495));
 assign mul_22_25_n_1471 = ((mul_22_25_n_1491 & mul_22_25_n_1492) | (mul_22_25_n_1490 & (mul_22_25_n_1491
    ^ mul_22_25_n_1492)));
 assign mul_22_25_n_1486 = (mul_22_25_n_1490 ^ (mul_22_25_n_1491 ^ mul_22_25_n_1492));
 assign mul_22_25_n_1468 = ((mul_22_25_n_1488 & mul_22_25_n_1489) | (mul_22_25_n_1487 & (mul_22_25_n_1488
    ^ mul_22_25_n_1489)));
 assign mul_22_25_n_1485 = (mul_22_25_n_1487 ^ (mul_22_25_n_1488 ^ mul_22_25_n_1489));
 assign mul_22_25_n_1804 = ((n_140 & n_88) | (n_143 & (n_140 ^ n_88)));
 assign mul_22_25_n_1768 = (n_143 ^ (n_140 ^ n_88));
 assign mul_22_25_n_1466 = ((mul_22_25_n_741 & mul_22_25_n_725) | (mul_22_25_n_752 & (mul_22_25_n_741
    ^ mul_22_25_n_725)));
 assign mul_22_25_n_1480 = (mul_22_25_n_752 ^ (mul_22_25_n_741 ^ mul_22_25_n_725));
 assign mul_22_25_n_1465 = ((mul_22_25_n_748 & mul_22_25_n_749) | (mul_22_25_n_502 & (mul_22_25_n_748
    ^ mul_22_25_n_749)));
 assign mul_22_25_n_1479 = (mul_22_25_n_502 ^ (mul_22_25_n_748 ^ mul_22_25_n_749));
 assign mul_22_25_n_1467 = ((mul_22_25_n_745 & mul_22_25_n_746) | (mul_22_25_n_744 & (mul_22_25_n_745
    ^ mul_22_25_n_746)));
 assign mul_22_25_n_1478 = (mul_22_25_n_744 ^ (mul_22_25_n_745 ^ mul_22_25_n_746));
 assign mul_22_25_n_1461 = ((mul_22_25_n_875 & mul_22_25_n_907) | (mul_22_25_n_1483 & (mul_22_25_n_875
    ^ mul_22_25_n_907)));
 assign mul_22_25_n_1476 = (mul_22_25_n_1483 ^ (mul_22_25_n_875 ^ mul_22_25_n_907));
 assign mul_22_25_n_1459 = ((mul_22_25_n_1481 & mul_22_25_n_1482) | (mul_22_25_n_1480 & (mul_22_25_n_1481
    ^ mul_22_25_n_1482)));
 assign mul_22_25_n_1474 = (mul_22_25_n_1480 ^ (mul_22_25_n_1481 ^ mul_22_25_n_1482));
 assign mul_22_25_n_1456 = ((mul_22_25_n_1478 & mul_22_25_n_1479) | (mul_22_25_n_1477 & (mul_22_25_n_1478
    ^ mul_22_25_n_1479)));
 assign mul_22_25_n_1473 = (mul_22_25_n_1477 ^ (mul_22_25_n_1478 ^ mul_22_25_n_1479));
 assign mul_22_25_n_1455 = ((mul_22_25_n_1475 & mul_22_25_n_1476) | (mul_22_25_n_1474 & (mul_22_25_n_1475
    ^ mul_22_25_n_1476)));
 assign mul_22_25_n_1470 = (mul_22_25_n_1474 ^ (mul_22_25_n_1475 ^ mul_22_25_n_1476));
 assign mul_22_25_n_1452 = ((mul_22_25_n_1472 & mul_22_25_n_1473) | (mul_22_25_n_1471 & (mul_22_25_n_1472
    ^ mul_22_25_n_1473)));
 assign mul_22_25_n_1469 = (mul_22_25_n_1471 ^ (mul_22_25_n_1472 ^ mul_22_25_n_1473));
 assign mul_22_25_n_1805 = ((n_136 & n_117) | (n_141 & (n_136 ^ n_117)));
 assign mul_22_25_n_1769 = (n_141 ^ (n_136 ^ n_117));
 assign mul_22_25_n_1449 = ((mul_22_25_n_665 & mul_22_25_n_723) | (mul_22_25_n_806 & (mul_22_25_n_665
    ^ mul_22_25_n_723)));
 assign mul_22_25_n_1464 = (mul_22_25_n_806 ^ (mul_22_25_n_665 ^ mul_22_25_n_723));
 assign mul_22_25_n_1450 = ((mul_22_25_n_731 & mul_22_25_n_732) | (mul_22_25_n_498 & (mul_22_25_n_731
    ^ mul_22_25_n_732)));
 assign mul_22_25_n_1463 = (mul_22_25_n_498 ^ (mul_22_25_n_731 ^ mul_22_25_n_732));
 assign mul_22_25_n_1451 = ((mul_22_25_n_639 & mul_22_25_n_729) | (mul_22_25_n_823 & (mul_22_25_n_639
    ^ mul_22_25_n_729)));
 assign mul_22_25_n_1462 = (mul_22_25_n_823 ^ (mul_22_25_n_639 ^ mul_22_25_n_729));
 assign mul_22_25_n_1445 = ((mul_22_25_n_874 & mul_22_25_n_906) | (mul_22_25_n_1467 & (mul_22_25_n_874
    ^ mul_22_25_n_906)));
 assign mul_22_25_n_1460 = (mul_22_25_n_1467 ^ (mul_22_25_n_874 ^ mul_22_25_n_906));
 assign mul_22_25_n_1444 = ((mul_22_25_n_1465 & mul_22_25_n_1466) | (mul_22_25_n_1464 & (mul_22_25_n_1465
    ^ mul_22_25_n_1466)));
 assign mul_22_25_n_1458 = (mul_22_25_n_1464 ^ (mul_22_25_n_1465 ^ mul_22_25_n_1466));
 assign mul_22_25_n_1441 = ((mul_22_25_n_1462 & mul_22_25_n_1463) | (mul_22_25_n_1461 & (mul_22_25_n_1462
    ^ mul_22_25_n_1463)));
 assign mul_22_25_n_1457 = (mul_22_25_n_1461 ^ (mul_22_25_n_1462 ^ mul_22_25_n_1463));
 assign mul_22_25_n_1439 = ((mul_22_25_n_1459 & mul_22_25_n_1460) | (mul_22_25_n_1458 & (mul_22_25_n_1459
    ^ mul_22_25_n_1460)));
 assign mul_22_25_n_1454 = (mul_22_25_n_1458 ^ (mul_22_25_n_1459 ^ mul_22_25_n_1460));
 assign mul_22_25_n_1436 = ((mul_22_25_n_1456 & mul_22_25_n_1457) | (mul_22_25_n_1455 & (mul_22_25_n_1456
    ^ mul_22_25_n_1457)));
 assign mul_22_25_n_1453 = (mul_22_25_n_1455 ^ (mul_22_25_n_1456 ^ mul_22_25_n_1457));
 assign mul_22_25_n_1806 = ((n_59 & n_55) | (n_137 & (n_59 ^ n_55)));
 assign mul_22_25_n_1770 = (n_137 ^ (n_59 ^ n_55));
 assign mul_22_25_n_1434 = ((mul_22_25_n_716 & mul_22_25_n_717) | (mul_22_25_n_677 & (mul_22_25_n_716
    ^ mul_22_25_n_717)));
 assign mul_22_25_n_1447 = (mul_22_25_n_677 ^ (mul_22_25_n_716 ^ mul_22_25_n_717));
 assign mul_22_25_n_1433 = ((mul_22_25_n_496 & mul_22_25_n_704) | (mul_22_25_n_1 & (mul_22_25_n_496 ^
    mul_22_25_n_704)));
 assign mul_22_25_n_1446 = (mul_22_25_n_1 ^ (mul_22_25_n_496 ^ mul_22_25_n_704));
 assign mul_22_25_n_1435 = ((mul_22_25_n_712 & mul_22_25_n_713) | (mul_22_25_n_721 & (mul_22_25_n_712
    ^ mul_22_25_n_713)));
 assign mul_22_25_n_1448 = (mul_22_25_n_721 ^ (mul_22_25_n_712 ^ mul_22_25_n_713));
 assign mul_22_25_n_1429 = ((mul_22_25_n_1451 & mul_22_25_n_868) | (mul_22_25_n_1450 & (mul_22_25_n_1451
    ^ mul_22_25_n_868)));
 assign mul_22_25_n_1443 = (mul_22_25_n_1450 ^ (mul_22_25_n_1451 ^ mul_22_25_n_868));
 assign mul_22_25_n_1428 = ((mul_22_25_n_1448 & mul_22_25_n_1449) | (mul_22_25_n_1447 & (mul_22_25_n_1448
    ^ mul_22_25_n_1449)));
 assign mul_22_25_n_1442 = (mul_22_25_n_1447 ^ (mul_22_25_n_1448 ^ mul_22_25_n_1449));
 assign mul_22_25_n_1424 = ((mul_22_25_n_910 & mul_22_25_n_1446) | (mul_22_25_n_1445 & (mul_22_25_n_910
    ^ mul_22_25_n_1446)));
 assign mul_22_25_n_1440 = (mul_22_25_n_1445 ^ (mul_22_25_n_910 ^ mul_22_25_n_1446));
 assign mul_22_25_n_1423 = ((mul_22_25_n_1443 & mul_22_25_n_1444) | (mul_22_25_n_1442 & (mul_22_25_n_1443
    ^ mul_22_25_n_1444)));
 assign mul_22_25_n_1438 = (mul_22_25_n_1442 ^ (mul_22_25_n_1443 ^ mul_22_25_n_1444));
 assign mul_22_25_n_1421 = ((mul_22_25_n_1440 & mul_22_25_n_1441) | (mul_22_25_n_1439 & (mul_22_25_n_1440
    ^ mul_22_25_n_1441)));
 assign mul_22_25_n_1437 = (mul_22_25_n_1439 ^ (mul_22_25_n_1440 ^ mul_22_25_n_1441));
 assign mul_22_25_n_1807 = ((n_46 & n_73) | (n_60 & (n_46 ^ n_73)));
 assign mul_22_25_n_1771 = (n_60 ^ (n_46 ^ n_73));
 assign mul_22_25_n_1419 = ((mul_22_25_n_787 & mul_22_25_n_755) | (mul_22_25_n_788 & (mul_22_25_n_787
    ^ mul_22_25_n_755)));
 assign mul_22_25_n_1432 = (mul_22_25_n_788 ^ (mul_22_25_n_787 ^ mul_22_25_n_755));
 assign mul_22_25_n_1418 = ((mul_22_25_n_497 & mul_22_25_n_812) | (mul_22_25_n_814 & (mul_22_25_n_497
    ^ mul_22_25_n_812)));
 assign mul_22_25_n_1431 = (mul_22_25_n_814 ^ (mul_22_25_n_497 ^ mul_22_25_n_812));
 assign mul_22_25_n_1417 = ((mul_22_25_n_818 & mul_22_25_n_615) | (mul_22_25_n_650 & (mul_22_25_n_818
    ^ mul_22_25_n_615)));
 assign mul_22_25_n_1430 = (mul_22_25_n_650 ^ (mul_22_25_n_818 ^ mul_22_25_n_615));
 assign mul_22_25_n_1412 = ((mul_22_25_n_1435 & mul_22_25_n_866) | (mul_22_25_n_878 & (mul_22_25_n_1435
    ^ mul_22_25_n_866)));
 assign mul_22_25_n_1426 = (mul_22_25_n_878 ^ (mul_22_25_n_1435 ^ mul_22_25_n_866));
 assign mul_22_25_n_1411 = ((mul_22_25_n_1433 & mul_22_25_n_1434) | (mul_22_25_n_1432 & (mul_22_25_n_1433
    ^ mul_22_25_n_1434)));
 assign mul_22_25_n_1427 = (mul_22_25_n_1432 ^ (mul_22_25_n_1433 ^ mul_22_25_n_1434));
 assign mul_22_25_n_1408 = ((mul_22_25_n_1430 & mul_22_25_n_1431) | (mul_22_25_n_1429 & (mul_22_25_n_1430
    ^ mul_22_25_n_1431)));
 assign mul_22_25_n_1425 = (mul_22_25_n_1429 ^ (mul_22_25_n_1430 ^ mul_22_25_n_1431));
 assign mul_22_25_n_1407 = ((mul_22_25_n_1427 & mul_22_25_n_1428) | (mul_22_25_n_1426 & (mul_22_25_n_1427
    ^ mul_22_25_n_1428)));
 assign mul_22_25_n_1422 = (mul_22_25_n_1426 ^ (mul_22_25_n_1427 ^ mul_22_25_n_1428));
 assign mul_22_25_n_1404 = ((mul_22_25_n_1424 & mul_22_25_n_1425) | (mul_22_25_n_1423 & (mul_22_25_n_1424
    ^ mul_22_25_n_1425)));
 assign mul_22_25_n_1420 = (mul_22_25_n_1423 ^ (mul_22_25_n_1424 ^ mul_22_25_n_1425));
 assign mul_22_25_n_1808 = ((n_47 & n_91) | (n_81 & (n_47 ^ n_91)));
 assign mul_22_25_n_1772 = (n_81 ^ (n_47 ^ n_91));
 assign mul_22_25_n_1403 = ((mul_22_25_n_754 & mul_22_25_n_6) | (mul_22_25_n_824 & (mul_22_25_n_754 ^
    mul_22_25_n_6)));
 assign mul_22_25_n_1415 = (mul_22_25_n_824 ^ (mul_22_25_n_754 ^ mul_22_25_n_6));
 assign mul_22_25_n_1402 = ((mul_22_25_n_651 & mul_22_25_n_825) | (mul_22_25_n_738 & (mul_22_25_n_651
    ^ mul_22_25_n_825)));
 assign mul_22_25_n_1414 = (mul_22_25_n_738 ^ (mul_22_25_n_651 ^ mul_22_25_n_825));
 assign mul_22_25_n_1401 = ((mul_22_25_n_827 & mul_22_25_n_463) | (mul_22_25_n_829 & (mul_22_25_n_827
    ^ mul_22_25_n_463)));
 assign mul_22_25_n_1416 = (mul_22_25_n_829 ^ (mul_22_25_n_827 ^ mul_22_25_n_463));
 assign mul_22_25_n_1397 = ((mul_22_25_n_865 & mul_22_25_n_676) | (mul_22_25_n_1419 & (mul_22_25_n_865
    ^ mul_22_25_n_676)));
 assign mul_22_25_n_1413 = (mul_22_25_n_1419 ^ (mul_22_25_n_865 ^ mul_22_25_n_676));
 assign mul_22_25_n_1396 = ((mul_22_25_n_1417 & mul_22_25_n_1418) | (mul_22_25_n_1416 & (mul_22_25_n_1417
    ^ mul_22_25_n_1418)));
 assign mul_22_25_n_1410 = (mul_22_25_n_1416 ^ (mul_22_25_n_1417 ^ mul_22_25_n_1418));
 assign mul_22_25_n_1393 = ((mul_22_25_n_1414 & mul_22_25_n_1415) | (mul_22_25_n_1413 & (mul_22_25_n_1414
    ^ mul_22_25_n_1415)));
 assign mul_22_25_n_1409 = (mul_22_25_n_1413 ^ (mul_22_25_n_1414 ^ mul_22_25_n_1415));
 assign mul_22_25_n_1392 = ((mul_22_25_n_1411 & mul_22_25_n_1412) | (mul_22_25_n_1410 & (mul_22_25_n_1411
    ^ mul_22_25_n_1412)));
 assign mul_22_25_n_1406 = (mul_22_25_n_1410 ^ (mul_22_25_n_1411 ^ mul_22_25_n_1412));
 assign mul_22_25_n_1389 = ((mul_22_25_n_1408 & mul_22_25_n_1409) | (mul_22_25_n_1407 & (mul_22_25_n_1408
    ^ mul_22_25_n_1409)));
 assign mul_22_25_n_1405 = (mul_22_25_n_1407 ^ (mul_22_25_n_1408 ^ mul_22_25_n_1409));
 assign mul_22_25_n_1809 = ((n_89 & n_87) | (n_82 & (n_89 ^ n_87)));
 assign mul_22_25_n_1773 = (n_82 ^ (n_89 ^ n_87));
 assign mul_22_25_n_1388 = ((mul_22_25_n_697 & mul_22_25_n_614) | (mul_22_25_n_467 & (mul_22_25_n_697
    ^ mul_22_25_n_614)));
 assign mul_22_25_n_1400 = (mul_22_25_n_467 ^ (mul_22_25_n_697 ^ mul_22_25_n_614));
 assign mul_22_25_n_1387 = ((mul_22_25_n_695 & mul_22_25_n_635) | (mul_22_25_n_693 & (mul_22_25_n_695
    ^ mul_22_25_n_635)));
 assign mul_22_25_n_1399 = (mul_22_25_n_693 ^ (mul_22_25_n_695 ^ mul_22_25_n_635));
 assign mul_22_25_n_1383 = ((mul_22_25_n_692 & mul_22_25_n_701) | (mul_22_25_n_0 & (mul_22_25_n_692 ^
    mul_22_25_n_701)));
 assign mul_22_25_n_1398 = (mul_22_25_n_0 ^ (mul_22_25_n_692 ^ mul_22_25_n_701));
 assign mul_22_25_n_1382 = ((mul_22_25_n_1402 & mul_22_25_n_1403) | (mul_22_25_n_1401 & (mul_22_25_n_1402
    ^ mul_22_25_n_1403)));
 assign mul_22_25_n_1395 = (mul_22_25_n_1401 ^ (mul_22_25_n_1402 ^ mul_22_25_n_1403));
 assign mul_22_25_n_1379 = ((mul_22_25_n_1399 & mul_22_25_n_1400) | (mul_22_25_n_1398 & (mul_22_25_n_1399
    ^ mul_22_25_n_1400)));
 assign mul_22_25_n_1394 = (mul_22_25_n_1398 ^ (mul_22_25_n_1399 ^ mul_22_25_n_1400));
 assign mul_22_25_n_1378 = ((mul_22_25_n_1396 & mul_22_25_n_1397) | (mul_22_25_n_1395 & (mul_22_25_n_1396
    ^ mul_22_25_n_1397)));
 assign mul_22_25_n_1391 = (mul_22_25_n_1395 ^ (mul_22_25_n_1396 ^ mul_22_25_n_1397));
 assign mul_22_25_n_1375 = ((mul_22_25_n_1393 & mul_22_25_n_1394) | (mul_22_25_n_1392 & (mul_22_25_n_1393
    ^ mul_22_25_n_1394)));
 assign mul_22_25_n_1390 = (mul_22_25_n_1392 ^ (mul_22_25_n_1393 ^ mul_22_25_n_1394));
 assign mul_22_25_n_1810 = ((n_129 & n_80) | (n_90 & (n_129 ^ n_80)));
 assign mul_22_25_n_1774 = (n_90 ^ (n_129 ^ n_80));
 assign mul_22_25_n_1374 = ((mul_22_25_n_685 & mul_22_25_n_811) | (mul_22_25_n_758 & (mul_22_25_n_685
    ^ mul_22_25_n_811)));
 assign mul_22_25_n_1386 = (mul_22_25_n_758 ^ (mul_22_25_n_685 ^ mul_22_25_n_811));
 assign mul_22_25_n_1373 = ((mul_22_25_n_475 & mul_22_25_n_683) | (mul_22_25_n_681 & (mul_22_25_n_475
    ^ mul_22_25_n_683)));
 assign mul_22_25_n_1384 = (mul_22_25_n_681 ^ (mul_22_25_n_475 ^ mul_22_25_n_683));
 assign mul_22_25_n_1372 = ((mul_22_25_n_680 & mul_22_25_n_652) | (mul_22_25_n_663 & (mul_22_25_n_680
    ^ mul_22_25_n_652)));
 assign mul_22_25_n_1385 = (mul_22_25_n_663 ^ (mul_22_25_n_680 ^ mul_22_25_n_652));
 assign mul_22_25_n_1368 = ((mul_22_25_n_1388 & mul_22_25_n_859) | (mul_22_25_n_1387 & (mul_22_25_n_1388
    ^ mul_22_25_n_859)));
 assign mul_22_25_n_1381 = (mul_22_25_n_1387 ^ (mul_22_25_n_1388 ^ mul_22_25_n_859));
 assign mul_22_25_n_1366 = ((mul_22_25_n_1385 & mul_22_25_n_1386) | (mul_22_25_n_1384 & (mul_22_25_n_1385
    ^ mul_22_25_n_1386)));
 assign mul_22_25_n_1380 = (mul_22_25_n_1384 ^ (mul_22_25_n_1385 ^ mul_22_25_n_1386));
 assign mul_22_25_n_1364 = ((mul_22_25_n_1382 & mul_22_25_n_1383) | (mul_22_25_n_1381 & (mul_22_25_n_1382
    ^ mul_22_25_n_1383)));
 assign mul_22_25_n_1377 = (mul_22_25_n_1381 ^ (mul_22_25_n_1382 ^ mul_22_25_n_1383));
 assign mul_22_25_n_1362 = ((mul_22_25_n_1379 & mul_22_25_n_1380) | (mul_22_25_n_1378 & (mul_22_25_n_1379
    ^ mul_22_25_n_1380)));
 assign mul_22_25_n_1376 = (mul_22_25_n_1378 ^ (mul_22_25_n_1379 ^ mul_22_25_n_1380));
 assign mul_22_25_n_1811 = ((n_106 & n_104) | (n_130 & (n_106 ^ n_104)));
 assign mul_22_25_n_1775 = (n_130 ^ (n_106 ^ n_104));
 assign mul_22_25_n_1360 = ((mul_22_25_n_470 & mul_22_25_n_673) | (mul_22_25_n_664 & (mul_22_25_n_470
    ^ mul_22_25_n_673)));
 assign mul_22_25_n_1370 = (mul_22_25_n_664 ^ (mul_22_25_n_470 ^ mul_22_25_n_673));
 assign mul_22_25_n_1361 = ((mul_22_25_n_668 & mul_22_25_n_669) | (mul_22_25_n_736 & (mul_22_25_n_668
    ^ mul_22_25_n_669)));
 assign mul_22_25_n_1371 = (mul_22_25_n_736 ^ (mul_22_25_n_668 ^ mul_22_25_n_669));
 assign mul_22_25_n_1356 = ((mul_22_25_n_850 & mul_22_25_n_786) | (mul_22_25_n_1374 & (mul_22_25_n_850
    ^ mul_22_25_n_786)));
 assign mul_22_25_n_1369 = (mul_22_25_n_1374 ^ (mul_22_25_n_850 ^ mul_22_25_n_786));
 assign mul_22_25_n_1354 = ((mul_22_25_n_1372 & mul_22_25_n_1373) | (mul_22_25_n_1371 & (mul_22_25_n_1372
    ^ mul_22_25_n_1373)));
 assign mul_22_25_n_1367 = (mul_22_25_n_1371 ^ (mul_22_25_n_1372 ^ mul_22_25_n_1373));
 assign mul_22_25_n_1353 = ((mul_22_25_n_1369 & mul_22_25_n_1370) | (mul_22_25_n_1368 & (mul_22_25_n_1369
    ^ mul_22_25_n_1370)));
 assign mul_22_25_n_1365 = (mul_22_25_n_1368 ^ (mul_22_25_n_1369 ^ mul_22_25_n_1370));
 assign mul_22_25_n_1350 = ((mul_22_25_n_1366 & mul_22_25_n_1367) | (mul_22_25_n_1365 & (mul_22_25_n_1366
    ^ mul_22_25_n_1367)));
 assign mul_22_25_n_1363 = (mul_22_25_n_1365 ^ (mul_22_25_n_1366 ^ mul_22_25_n_1367));
 assign mul_22_25_n_1812 = ((n_148 & n_105) | (n_107 & (n_148 ^ n_105)));
 assign mul_22_25_n_1776 = (n_107 ^ (n_148 ^ n_105));
 assign mul_22_25_n_1349 = ((mul_22_25_n_670 & mul_22_25_n_813) | (mul_22_25_n_660 & (mul_22_25_n_670
    ^ mul_22_25_n_813)));
 assign mul_22_25_n_1359 = (mul_22_25_n_660 ^ (mul_22_25_n_670 ^ mul_22_25_n_813));
 assign mul_22_25_n_1348 = ((mul_22_25_n_659 & mul_22_25_n_471) | (mul_22_25_n_641 & (mul_22_25_n_659
    ^ mul_22_25_n_471)));
 assign mul_22_25_n_1358 = (mul_22_25_n_641 ^ (mul_22_25_n_659 ^ mul_22_25_n_471));
 assign mul_22_25_n_1345 = ((mul_22_25_n_618 & mul_22_25_n_791) | (mul_22_25_n_851 & (mul_22_25_n_618
    ^ mul_22_25_n_791)));
 assign mul_22_25_n_1357 = (mul_22_25_n_851 ^ (mul_22_25_n_618 ^ mul_22_25_n_791));
 assign mul_22_25_n_1343 = ((mul_22_25_n_1360 & mul_22_25_n_1361) | (mul_22_25_n_1359 & (mul_22_25_n_1360
    ^ mul_22_25_n_1361)));
 assign mul_22_25_n_1355 = (mul_22_25_n_1359 ^ (mul_22_25_n_1360 ^ mul_22_25_n_1361));
 assign mul_22_25_n_1341 = ((mul_22_25_n_1357 & mul_22_25_n_1358) | (mul_22_25_n_1356 & (mul_22_25_n_1357
    ^ mul_22_25_n_1358)));
 assign mul_22_25_n_1352 = (mul_22_25_n_1356 ^ (mul_22_25_n_1357 ^ mul_22_25_n_1358));
 assign mul_22_25_n_1339 = ((mul_22_25_n_1354 & mul_22_25_n_1355) | (mul_22_25_n_1353 & (mul_22_25_n_1354
    ^ mul_22_25_n_1355)));
 assign mul_22_25_n_1351 = (mul_22_25_n_1353 ^ (mul_22_25_n_1354 ^ mul_22_25_n_1355));
 assign mul_22_25_n_1778 = ((n_147 & n_151) | (n_149 & (n_147 ^ n_151)));
 assign mul_22_25_n_1777 = (n_149 ^ (n_147 ^ n_151));
 assign mul_22_25_n_1338 = ((mul_22_25_n_634 & mul_22_25_n_637) | (mul_22_25_n_702 & (mul_22_25_n_634
    ^ mul_22_25_n_637)));
 assign mul_22_25_n_1346 = (mul_22_25_n_702 ^ (mul_22_25_n_634 ^ mul_22_25_n_637));
 assign mul_22_25_n_1337 = ((mul_22_25_n_699 & mul_22_25_n_657) | (mul_22_25_n_465 & (mul_22_25_n_699
    ^ mul_22_25_n_657)));
 assign mul_22_25_n_1347 = (mul_22_25_n_465 ^ (mul_22_25_n_699 ^ mul_22_25_n_657));
 assign mul_22_25_n_1333 = ((mul_22_25_n_1349 & mul_22_25_n_861) | (mul_22_25_n_1348 & (mul_22_25_n_1349
    ^ mul_22_25_n_861)));
 assign mul_22_25_n_1344 = (mul_22_25_n_1348 ^ (mul_22_25_n_1349 ^ mul_22_25_n_861));
 assign mul_22_25_n_1332 = ((mul_22_25_n_1346 & mul_22_25_n_1347) | (mul_22_25_n_1345 & (mul_22_25_n_1346
    ^ mul_22_25_n_1347)));
 assign mul_22_25_n_1342 = (mul_22_25_n_1345 ^ (mul_22_25_n_1346 ^ mul_22_25_n_1347));
 assign mul_22_25_n_1329 = ((mul_22_25_n_1343 & mul_22_25_n_1344) | (mul_22_25_n_1342 & (mul_22_25_n_1343
    ^ mul_22_25_n_1344)));
 assign mul_22_25_n_1340 = (mul_22_25_n_1342 ^ (mul_22_25_n_1343 ^ mul_22_25_n_1344));
 assign mul_22_25_n_1814 = ((mul_22_25_n_1340 & mul_22_25_n_1341) | (mul_22_25_n_1339 & (mul_22_25_n_1340
    ^ mul_22_25_n_1341)));
 assign mul_22_25_n_1813 = (mul_22_25_n_1339 ^ (mul_22_25_n_1340 ^ mul_22_25_n_1341));
 assign mul_22_25_n_1327 = ((mul_22_25_n_580 & mul_22_25_n_805) | (mul_22_25_n_604 & (mul_22_25_n_580
    ^ mul_22_25_n_805)));
 assign mul_22_25_n_1335 = (mul_22_25_n_604 ^ (mul_22_25_n_580 ^ mul_22_25_n_805));
 assign mul_22_25_n_1328 = ((mul_22_25_n_671 & mul_22_25_n_648) | (mul_22_25_n_679 & (mul_22_25_n_671
    ^ mul_22_25_n_648)));
 assign mul_22_25_n_1336 = (mul_22_25_n_679 ^ (mul_22_25_n_671 ^ mul_22_25_n_648));
 assign mul_22_25_n_1324 = ((mul_22_25_n_860 & mul_22_25_n_459) | (mul_22_25_n_1338 & (mul_22_25_n_860
    ^ mul_22_25_n_459)));
 assign mul_22_25_n_1334 = (mul_22_25_n_1338 ^ (mul_22_25_n_860 ^ mul_22_25_n_459));
 assign mul_22_25_n_1323 = ((mul_22_25_n_1336 & mul_22_25_n_1337) | (mul_22_25_n_1335 & (mul_22_25_n_1336
    ^ mul_22_25_n_1337)));
 assign mul_22_25_n_1331 = (mul_22_25_n_1335 ^ (mul_22_25_n_1336 ^ mul_22_25_n_1337));
 assign mul_22_25_n_1320 = ((mul_22_25_n_1333 & mul_22_25_n_1334) | (mul_22_25_n_1332 & (mul_22_25_n_1333
    ^ mul_22_25_n_1334)));
 assign mul_22_25_n_1330 = (mul_22_25_n_1332 ^ (mul_22_25_n_1333 ^ mul_22_25_n_1334));
 assign mul_22_25_n_1815 = ((mul_22_25_n_1330 & mul_22_25_n_1331) | (mul_22_25_n_1329 & (mul_22_25_n_1330
    ^ mul_22_25_n_1331)));
 assign mul_22_25_n_1779 = (mul_22_25_n_1329 ^ (mul_22_25_n_1330 ^ mul_22_25_n_1331));
 assign mul_22_25_n_1319 = ((mul_22_25_n_599 & mul_22_25_n_563) | (mul_22_25_n_808 & (mul_22_25_n_599
    ^ mul_22_25_n_563)));
 assign mul_22_25_n_1326 = (mul_22_25_n_808 ^ (mul_22_25_n_599 ^ mul_22_25_n_563));
 assign mul_22_25_n_1316 = ((mul_22_25_n_640 & mul_22_25_n_500) | (mul_22_25_n_862 & (mul_22_25_n_640
    ^ mul_22_25_n_500)));
 assign mul_22_25_n_1325 = (mul_22_25_n_862 ^ (mul_22_25_n_640 ^ mul_22_25_n_500));
 assign mul_22_25_n_1314 = ((mul_22_25_n_1327 & mul_22_25_n_1328) | (mul_22_25_n_1326 & (mul_22_25_n_1327
    ^ mul_22_25_n_1328)));
 assign mul_22_25_n_1322 = (mul_22_25_n_1326 ^ (mul_22_25_n_1327 ^ mul_22_25_n_1328));
 assign mul_22_25_n_1312 = ((mul_22_25_n_1324 & mul_22_25_n_1325) | (mul_22_25_n_1323 & (mul_22_25_n_1324
    ^ mul_22_25_n_1325)));
 assign mul_22_25_n_1321 = (mul_22_25_n_1323 ^ (mul_22_25_n_1324 ^ mul_22_25_n_1325));
 assign mul_22_25_n_1816 = ((mul_22_25_n_1321 & mul_22_25_n_1322) | (mul_22_25_n_1320 & (mul_22_25_n_1321
    ^ mul_22_25_n_1322)));
 assign mul_22_25_n_1780 = (mul_22_25_n_1320 ^ (mul_22_25_n_1321 ^ mul_22_25_n_1322));
 assign mul_22_25_n_1310 = ((mul_22_25_n_763 & mul_22_25_n_815) | (mul_22_25_n_753 & (mul_22_25_n_763
    ^ mul_22_25_n_815)));
 assign mul_22_25_n_1317 = (mul_22_25_n_753 ^ (mul_22_25_n_763 ^ mul_22_25_n_815));
 assign mul_22_25_n_1311 = ((mul_22_25_n_569 & mul_22_25_n_645) | (mul_22_25_n_464 & (mul_22_25_n_569
    ^ mul_22_25_n_645)));
 assign mul_22_25_n_1318 = (mul_22_25_n_464 ^ (mul_22_25_n_569 ^ mul_22_25_n_645));
 assign mul_22_25_n_1307 = ((mul_22_25_n_1319 & mul_22_25_n_863) | (mul_22_25_n_1318 & (mul_22_25_n_1319
    ^ mul_22_25_n_863)));
 assign mul_22_25_n_1315 = (mul_22_25_n_1318 ^ (mul_22_25_n_1319 ^ mul_22_25_n_863));
 assign mul_22_25_n_1305 = ((mul_22_25_n_1316 & mul_22_25_n_1317) | (mul_22_25_n_1315 & (mul_22_25_n_1316
    ^ mul_22_25_n_1317)));
 assign mul_22_25_n_1313 = (mul_22_25_n_1315 ^ (mul_22_25_n_1316 ^ mul_22_25_n_1317));
 assign mul_22_25_n_1817 = ((mul_22_25_n_1313 & mul_22_25_n_1314) | (mul_22_25_n_1312 & (mul_22_25_n_1313
    ^ mul_22_25_n_1314)));
 assign mul_22_25_n_1781 = (mul_22_25_n_1312 ^ (mul_22_25_n_1313 ^ mul_22_25_n_1314));
 assign mul_22_25_n_1304 = ((mul_22_25_n_462 & mul_22_25_n_631) | (mul_22_25_n_810 & (mul_22_25_n_462
    ^ mul_22_25_n_631)));
 assign mul_22_25_n_1309 = (mul_22_25_n_810 ^ (mul_22_25_n_462 ^ mul_22_25_n_631));
 assign mul_22_25_n_1301 = ((mul_22_25_n_856 & mul_22_25_n_629) | (mul_22_25_n_1311 & (mul_22_25_n_856
    ^ mul_22_25_n_629)));
 assign mul_22_25_n_1308 = (mul_22_25_n_1311 ^ (mul_22_25_n_856 ^ mul_22_25_n_629));
 assign mul_22_25_n_1299 = ((mul_22_25_n_1309 & mul_22_25_n_1310) | (mul_22_25_n_1308 & (mul_22_25_n_1309
    ^ mul_22_25_n_1310)));
 assign mul_22_25_n_1306 = (mul_22_25_n_1308 ^ (mul_22_25_n_1309 ^ mul_22_25_n_1310));
 assign mul_22_25_n_1783 = ((mul_22_25_n_1306 & mul_22_25_n_1307) | (mul_22_25_n_1305 & (mul_22_25_n_1306
    ^ mul_22_25_n_1307)));
 assign mul_22_25_n_1782 = (mul_22_25_n_1305 ^ (mul_22_25_n_1306 ^ mul_22_25_n_1307));
 assign mul_22_25_n_1298 = ((mul_22_25_n_623 & mul_22_25_n_7) | (mul_22_25_n_624 & (mul_22_25_n_623 ^
    mul_22_25_n_7)));
 assign mul_22_25_n_1303 = (mul_22_25_n_624 ^ (mul_22_25_n_623 ^ mul_22_25_n_7));
 assign mul_22_25_n_1296 = ((mul_22_25_n_636 & mul_22_25_n_474) | (mul_22_25_n_857 & (mul_22_25_n_636
    ^ mul_22_25_n_474)));
 assign mul_22_25_n_1302 = (mul_22_25_n_857 ^ (mul_22_25_n_636 ^ mul_22_25_n_474));
 assign mul_22_25_n_1294 = ((mul_22_25_n_1303 & mul_22_25_n_1304) | (mul_22_25_n_1302 & (mul_22_25_n_1303
    ^ mul_22_25_n_1304)));
 assign mul_22_25_n_1300 = (mul_22_25_n_1302 ^ (mul_22_25_n_1303 ^ mul_22_25_n_1304));
 assign mul_22_25_n_1784 = ((mul_22_25_n_1300 & mul_22_25_n_1301) | (mul_22_25_n_1299 & (mul_22_25_n_1300
    ^ mul_22_25_n_1301)));
 assign mul_22_25_n_1265 = (mul_22_25_n_1299 ^ (mul_22_25_n_1300 ^ mul_22_25_n_1301));
 assign mul_22_25_n_1293 = ((mul_22_25_n_619 & mul_22_25_n_468) | (mul_22_25_n_632 & (mul_22_25_n_619
    ^ mul_22_25_n_468)));
 assign mul_22_25_n_1297 = (mul_22_25_n_632 ^ (mul_22_25_n_619 ^ mul_22_25_n_468));
 assign mul_22_25_n_1290 = ((mul_22_25_n_1298 & mul_22_25_n_854) | (mul_22_25_n_1297 & (mul_22_25_n_1298
    ^ mul_22_25_n_854)));
 assign mul_22_25_n_1295 = (mul_22_25_n_1297 ^ (mul_22_25_n_1298 ^ mul_22_25_n_854));
 assign mul_22_25_n_1270 = ((mul_22_25_n_1295 & mul_22_25_n_1296) | (mul_22_25_n_1294 & (mul_22_25_n_1295
    ^ mul_22_25_n_1296)));
 assign mul_22_25_n_1818 = (mul_22_25_n_1294 ^ (mul_22_25_n_1295 ^ mul_22_25_n_1296));
 assign mul_22_25_n_1289 = ((mul_22_25_n_773 & mul_22_25_n_809) | (mul_22_25_n_466 & (mul_22_25_n_773
    ^ mul_22_25_n_809)));
 assign mul_22_25_n_1292 = (mul_22_25_n_466 ^ (mul_22_25_n_773 ^ mul_22_25_n_809));
 assign mul_22_25_n_1287 = ((mul_22_25_n_855 & mul_22_25_n_581) | (mul_22_25_n_1293 & (mul_22_25_n_855
    ^ mul_22_25_n_581)));
 assign mul_22_25_n_1291 = (mul_22_25_n_1293 ^ (mul_22_25_n_855 ^ mul_22_25_n_581));
 assign mul_22_25_n_1269 = ((mul_22_25_n_1291 & mul_22_25_n_1292) | (mul_22_25_n_1290 & (mul_22_25_n_1291
    ^ mul_22_25_n_1292)));
 assign mul_22_25_n_1268 = (mul_22_25_n_1290 ^ (mul_22_25_n_1291 ^ mul_22_25_n_1292));
 assign mul_22_25_n_1285 = ((mul_22_25_n_472 & mul_22_25_n_767) | (mul_22_25_n_852 & (mul_22_25_n_472
    ^ mul_22_25_n_767)));
 assign mul_22_25_n_1288 = (mul_22_25_n_852 ^ (mul_22_25_n_472 ^ mul_22_25_n_767));
 assign mul_22_25_n_1267 = ((mul_22_25_n_1288 & mul_22_25_n_1289) | (mul_22_25_n_1287 & (mul_22_25_n_1288
    ^ mul_22_25_n_1289)));
 assign mul_22_25_n_1266 = (mul_22_25_n_1287 ^ (mul_22_25_n_1288 ^ mul_22_25_n_1289));
 assign mul_22_25_n_1284 = ((mul_22_25_n_586 & mul_22_25_n_807) | (mul_22_25_n_499 & (mul_22_25_n_586
    ^ mul_22_25_n_807)));
 assign mul_22_25_n_1286 = (mul_22_25_n_499 ^ (mul_22_25_n_586 ^ mul_22_25_n_807));
 assign mul_22_25_n_1275 = ((mul_22_25_n_1286 & mul_22_25_n_853) | (mul_22_25_n_1285 & (mul_22_25_n_1286
    ^ mul_22_25_n_853)));
 assign mul_22_25_n_1819 = (mul_22_25_n_1285 ^ (mul_22_25_n_1286 ^ mul_22_25_n_853));
 assign mul_22_25_n_19 = ~(n_114 | (~mul_22_25_n_1245 & n_115));
 assign asc001_47_ = (mul_22_25_n_969 ^ mul_22_25_n_1263);
 assign mul_22_25_n_1263 = ~(n_102 | (mul_22_25_n_1257 & n_103));
 assign asc001_46_ = ~(mul_22_25_n_968 ^ mul_22_25_n_1257);
 assign asc001_45_ = (mul_22_25_n_1020 ^ mul_22_25_n_19);
 assign asc001_43_ = (mul_22_25_n_1023 ^ mul_22_25_n_1255);
 assign asc001_39_ = (mul_22_25_n_1139 ^ mul_22_25_n_1254);
 assign asc001_49_ = (n_152 ^ mul_22_25_n_1233);
 assign asc001_44_ = (mul_22_25_n_1024 ^ mul_22_25_n_1245);
 assign mul_22_25_n_1255 = ~(n_43 | (mul_22_25_n_1246 & n_68));
 assign mul_22_25_n_1254 = ~(mul_22_25_n_1118 | (mul_22_25_n_1247 & mul_22_25_n_1112));
 assign mul_22_25_n_1257 = ~(mul_22_25_n_1039 & (mul_22_25_n_1245 | mul_22_25_n_1035));
 assign asc001_42_ = ~(mul_22_25_n_1022 ^ mul_22_25_n_1246);
 assign asc001_41_ = (mul_22_25_n_1021 ^ mul_22_25_n_1242);
 assign asc001_38_ = ~(mul_22_25_n_1138 ^ mul_22_25_n_1247);
 assign asc001_37_ = (mul_22_25_n_1137 ^ mul_22_25_n_1243);
 assign asc001_35_ = (mul_22_25_n_1135 ^ mul_22_25_n_1240);
 assign asc001_31_ = (mul_22_25_n_1140 ^ mul_22_25_n_1241);
 assign asc001_27_ = (mul_22_25_n_1148 ^ mul_22_25_n_1226);
 assign mul_22_25_n_1243 = ~(mul_22_25_n_1107 | (mul_22_25_n_1229 & mul_22_25_n_1101));
 assign mul_22_25_n_1242 = ~(n_144 | (mul_22_25_n_1228 & n_58));
 assign mul_22_25_n_1241 = ~(mul_22_25_n_1120 | (mul_22_25_n_1224 & mul_22_25_n_1116));
 assign mul_22_25_n_1240 = ~(mul_22_25_n_1098 | (mul_22_25_n_1231 & mul_22_25_n_1093));
 assign mul_22_25_n_1247 = ~(mul_22_25_n_1172 & (mul_22_25_n_1230 | mul_22_25_n_1159));
 assign mul_22_25_n_1246 = ~(mul_22_25_n_1171 & (mul_22_25_n_1227 | mul_22_25_n_1164));
 assign mul_22_25_n_1245 = ~(mul_22_25_n_1192 | (mul_22_25_n_1228 & mul_22_25_n_1173));
 assign asc001_30_ = ~(mul_22_25_n_1131 ^ mul_22_25_n_1224);
 assign asc001_36_ = ~((mul_22_25_n_1229 & ~mul_22_25_n_1136) | (mul_22_25_n_1230 & mul_22_25_n_1136));
 assign asc001_34_ = ~(mul_22_25_n_1134 ^ mul_22_25_n_1231);
 assign asc001_33_ = (mul_22_25_n_1133 ^ mul_22_25_n_1225);
 assign asc001_40_ = ~((mul_22_25_n_1228 & ~mul_22_25_n_1127) | (mul_22_25_n_1227 & mul_22_25_n_1127));
 assign asc001_29_ = (mul_22_25_n_1130 ^ mul_22_25_n_1218);
 assign mul_22_25_n_1233 = ~(n_139 | (mul_22_25_n_1232 & n_138));
 assign mul_22_25_n_1229 = ~mul_22_25_n_1230;
 assign mul_22_25_n_1227 = ~mul_22_25_n_1228;
 assign mul_22_25_n_1226 = ~(mul_22_25_n_1115 | (mul_22_25_n_1217 & mul_22_25_n_1113));
 assign mul_22_25_n_1225 = ~(mul_22_25_n_1091 | (mul_22_25_n_1210 & mul_22_25_n_1088));
 assign mul_22_25_n_1232 = ~(mul_22_25_n_1214 & (mul_22_25_n_1189 | (mul_22_25_n_1182 | mul_22_25_n_1211)));
 assign mul_22_25_n_1231 = ~(mul_22_25_n_1169 & (mul_22_25_n_1211 | mul_22_25_n_1145));
 assign mul_22_25_n_1230 = ~(mul_22_25_n_1191 | (mul_22_25_n_1210 & mul_22_25_n_1174));
 assign mul_22_25_n_1228 = ~(mul_22_25_n_1201 & (mul_22_25_n_1211 | mul_22_25_n_1182));
 assign asc001_28_ = (mul_22_25_n_1129 ^ mul_22_25_n_1213);
 assign asc001_32_ = ~((mul_22_25_n_1210 & ~mul_22_25_n_1132) | (mul_22_25_n_1211 & mul_22_25_n_1132));
 assign asc001_26_ = ~(mul_22_25_n_1155 ^ mul_22_25_n_1217);
 assign asc001_25_ = (mul_22_25_n_1154 ^ mul_22_25_n_1216);
 assign asc001_23_ = ~(mul_22_25_n_1152 ^ mul_22_25_n_1215);
 assign mul_22_25_n_1218 = ~(mul_22_25_n_1106 | (mul_22_25_n_1212 & mul_22_25_n_1117));
 assign mul_22_25_n_1224 = ~(mul_22_25_n_1179 & (mul_22_25_n_1213 | mul_22_25_n_1163));
 assign mul_22_25_n_1217 = ~(mul_22_25_n_1168 & (mul_22_25_n_1203 | mul_22_25_n_1160));
 assign mul_22_25_n_1216 = (~mul_22_25_n_1109 & (mul_22_25_n_1203 | mul_22_25_n_1087));
 assign mul_22_25_n_1215 = ~(mul_22_25_n_1100 & (mul_22_25_n_1202 | mul_22_25_n_1092));
 assign mul_22_25_n_1214 = ~(mul_22_25_n_1049 | (mul_22_25_n_1206 | (mul_22_25_n_1192 & mul_22_25_n_1041)));
 assign mul_22_25_n_1213 = ~mul_22_25_n_1212;
 assign mul_22_25_n_1212 = ~(mul_22_25_n_1193 & (mul_22_25_n_1203 | mul_22_25_n_1177));
 assign mul_22_25_n_1210 = ~mul_22_25_n_1211;
 assign mul_22_25_n_1211 = ~(mul_22_25_n_1205 | (mul_22_25_n_1195 & mul_22_25_n_1190));
 assign asc001_24_ = (mul_22_25_n_1153 ^ mul_22_25_n_1203);
 assign asc001_22_ = (mul_22_25_n_1151 ^ mul_22_25_n_1202);
 assign asc001_21_ = ~(mul_22_25_n_1150 ^ mul_22_25_n_1200);
 assign mul_22_25_n_1206 = ~(mul_22_25_n_1201 | mul_22_25_n_1189);
 assign mul_22_25_n_1205 = ~(mul_22_25_n_1194 & (mul_22_25_n_1204 & (mul_22_25_n_1193 | mul_22_25_n_1178)));
 assign mul_22_25_n_1204 = ~(mul_22_25_n_1198 & mul_22_25_n_1190);
 assign mul_22_25_n_1203 = ~(mul_22_25_n_1195 | mul_22_25_n_1198);
 assign mul_22_25_n_1202 = ~(mul_22_25_n_1170 | (mul_22_25_n_1196 & mul_22_25_n_1157));
 assign mul_22_25_n_1201 = ~(mul_22_25_n_1187 | (mul_22_25_n_1166 | (mul_22_25_n_1191 & mul_22_25_n_1176)));
 assign mul_22_25_n_1200 = ~(mul_22_25_n_1099 | (mul_22_25_n_1196 & mul_22_25_n_1097));
 assign asc001_20_ = ~(mul_22_25_n_1149 ^ mul_22_25_n_1196);
 assign mul_22_25_n_1198 = ~(mul_22_25_n_1185 & (mul_22_25_n_1167 & (mul_22_25_n_1184 | mul_22_25_n_1175)));
 assign asc001_19_ = ~(mul_22_25_n_1147 ^ mul_22_25_n_1180);
 assign mul_22_25_n_1196 = ~(mul_22_25_n_1183 & mul_22_25_n_1184);
 assign mul_22_25_n_1195 = ~(mul_22_25_n_1183 | mul_22_25_n_1175);
 assign mul_22_25_n_1194 = ~(mul_22_25_n_1123 | (mul_22_25_n_1186 | (mul_22_25_n_1110 & mul_22_25_n_1120)));
 assign mul_22_25_n_1193 = ~(mul_22_25_n_1126 | (mul_22_25_n_1188 | (mul_22_25_n_1114 & mul_22_25_n_1115)));
 assign mul_22_25_n_1192 = ~(mul_22_25_n_1034 & (n_110 & (mul_22_25_n_1171 | mul_22_25_n_1028)));
 assign mul_22_25_n_1191 = ~(mul_22_25_n_1156 & (mul_22_25_n_1104 & (mul_22_25_n_1169 | mul_22_25_n_1146)));
 assign mul_22_25_n_1188 = ~(mul_22_25_n_1168 | mul_22_25_n_1162);
 assign mul_22_25_n_1187 = ~(mul_22_25_n_1172 | mul_22_25_n_1161);
 assign mul_22_25_n_1186 = ~(mul_22_25_n_1179 | mul_22_25_n_1165);
 assign mul_22_25_n_1185 = ~(mul_22_25_n_1170 & mul_22_25_n_1158);
 assign mul_22_25_n_1190 = ~(mul_22_25_n_1178 | mul_22_25_n_1177);
 assign mul_22_25_n_1189 = ~(mul_22_25_n_1041 & mul_22_25_n_1173);
 assign asc001_17_ = ~(mul_22_25_n_1033 ^ mul_22_25_n_1128);
 assign mul_22_25_n_1184 = ~(mul_22_25_n_1142 | (mul_22_25_n_1105 | (mul_22_25_n_1040 & mul_22_25_n_1144)));
 assign mul_22_25_n_1183 = ~(mul_22_25_n_1144 & (mul_22_25_n_1027 & mul_22_25_n_1067));
 assign mul_22_25_n_1182 = ~(mul_22_25_n_1176 & mul_22_25_n_1174);
 assign mul_22_25_n_1180 = ~(mul_22_25_n_1046 & (mul_22_25_n_1143 | mul_22_25_n_1045));
 assign mul_22_25_n_1179 = ~(mul_22_25_n_1121 | (mul_22_25_n_1119 & mul_22_25_n_1106));
 assign mul_22_25_n_1178 = (mul_22_25_n_1165 | mul_22_25_n_1163);
 assign mul_22_25_n_1177 = (mul_22_25_n_1162 | mul_22_25_n_1160);
 assign mul_22_25_n_1176 = ~(mul_22_25_n_1161 | mul_22_25_n_1159);
 assign mul_22_25_n_1175 = ~(mul_22_25_n_1158 & mul_22_25_n_1157);
 assign mul_22_25_n_1174 = ~(mul_22_25_n_1146 | mul_22_25_n_1145);
 assign mul_22_25_n_1173 = ~(mul_22_25_n_1028 | mul_22_25_n_1164);
 assign mul_22_25_n_1167 = (~mul_22_25_n_15 & (mul_22_25_n_1095 | mul_22_25_n_1100));
 assign mul_22_25_n_1166 = (~mul_22_25_n_1122 | (mul_22_25_n_16 & mul_22_25_n_1118));
 assign mul_22_25_n_1172 = ~(mul_22_25_n_1125 | (mul_22_25_n_1096 & mul_22_25_n_1107));
 assign mul_22_25_n_1171 = ~(n_42 | (n_61 & n_144));
 assign mul_22_25_n_1170 = (~mul_22_25_n_1103 | (mul_22_25_n_14 & mul_22_25_n_1099));
 assign mul_22_25_n_1169 = ~(mul_22_25_n_1102 | (mul_22_25_n_1090 & mul_22_25_n_1091));
 assign mul_22_25_n_1168 = ~(mul_22_25_n_1124 | (mul_22_25_n_1108 & mul_22_25_n_1109));
 assign mul_22_25_n_1156 = ~(mul_22_25_n_13 & mul_22_25_n_1098);
 assign mul_22_25_n_1155 = ~(mul_22_25_n_1113 & ~mul_22_25_n_1115);
 assign mul_22_25_n_1154 = ~(mul_22_25_n_1108 & ~mul_22_25_n_1124);
 assign mul_22_25_n_1153 = (mul_22_25_n_1087 | mul_22_25_n_1109);
 assign mul_22_25_n_1152 = (mul_22_25_n_1095 | mul_22_25_n_15);
 assign mul_22_25_n_1151 = ~(mul_22_25_n_1100 & ~mul_22_25_n_1092);
 assign mul_22_25_n_1150 = (mul_22_25_n_14 & mul_22_25_n_1103);
 assign mul_22_25_n_1165 = ~(mul_22_25_n_1110 & mul_22_25_n_1116);
 assign mul_22_25_n_1149 = ~(~mul_22_25_n_1099 & mul_22_25_n_1097);
 assign mul_22_25_n_1148 = ~(mul_22_25_n_1114 & ~mul_22_25_n_1126);
 assign mul_22_25_n_1164 = ~(n_61 & n_58);
 assign mul_22_25_n_1163 = ~(mul_22_25_n_1119 & mul_22_25_n_1117);
 assign mul_22_25_n_1162 = ~(mul_22_25_n_1114 & mul_22_25_n_1113);
 assign mul_22_25_n_1161 = ~(mul_22_25_n_16 & mul_22_25_n_1112);
 assign mul_22_25_n_1160 = ~(mul_22_25_n_1108 & ~mul_22_25_n_1087);
 assign mul_22_25_n_1159 = ~(mul_22_25_n_1096 & mul_22_25_n_1101);
 assign mul_22_25_n_1158 = ~(mul_22_25_n_1095 | mul_22_25_n_1092);
 assign mul_22_25_n_1147 = ~(~mul_22_25_n_1105 & mul_22_25_n_1094);
 assign mul_22_25_n_1157 = (mul_22_25_n_14 & mul_22_25_n_1097);
 assign mul_22_25_n_1142 = ~(~mul_22_25_n_1094 | mul_22_25_n_1046);
 assign asc001_16_ = ~(mul_22_25_n_1032 ^ mul_22_25_n_1067);
 assign mul_22_25_n_1140 = ~(mul_22_25_n_1110 & ~mul_22_25_n_1123);
 assign mul_22_25_n_1139 = ~(mul_22_25_n_16 & mul_22_25_n_1122);
 assign mul_22_25_n_1138 = ~(~mul_22_25_n_1118 & mul_22_25_n_1112);
 assign mul_22_25_n_1137 = ~(mul_22_25_n_1096 & ~mul_22_25_n_1125);
 assign mul_22_25_n_1136 = ~(~mul_22_25_n_1107 & mul_22_25_n_1101);
 assign mul_22_25_n_1135 = ~(mul_22_25_n_13 & mul_22_25_n_1104);
 assign mul_22_25_n_1134 = ~(~mul_22_25_n_1098 & mul_22_25_n_1093);
 assign mul_22_25_n_1133 = ~(mul_22_25_n_1090 & ~mul_22_25_n_1102);
 assign mul_22_25_n_1132 = ~(~mul_22_25_n_1091 & mul_22_25_n_1088);
 assign mul_22_25_n_1146 = ~(mul_22_25_n_13 & mul_22_25_n_1093);
 assign mul_22_25_n_1145 = ~(mul_22_25_n_1090 & mul_22_25_n_1088);
 assign mul_22_25_n_1131 = ~(mul_22_25_n_1116 & ~mul_22_25_n_1120);
 assign mul_22_25_n_1130 = ~(mul_22_25_n_1119 & ~mul_22_25_n_1121);
 assign mul_22_25_n_1129 = ~(mul_22_25_n_1117 & ~mul_22_25_n_1106);
 assign mul_22_25_n_1144 = ~(~mul_22_25_n_1094 | mul_22_25_n_1045);
 assign mul_22_25_n_1128 = (~n_57 | (mul_22_25_n_1067 & n_95));
 assign mul_22_25_n_1127 = ~(~n_144 & n_58);
 assign mul_22_25_n_1143 = ~(mul_22_25_n_1040 | (mul_22_25_n_1067 & mul_22_25_n_1027));
 assign mul_22_25_n_1126 = ~(mul_22_25_n_1074 | mul_22_25_n_1075);
 assign mul_22_25_n_1125 = ~(mul_22_25_n_1065 | mul_22_25_n_1068);
 assign mul_22_25_n_1124 = ~(mul_22_25_n_1069 | mul_22_25_n_1070);
 assign mul_22_25_n_1123 = ~(mul_22_25_n_1083 | mul_22_25_n_1084);
 assign mul_22_25_n_1122 = ~(n_150 & mul_22_25_n_1778);
 assign mul_22_25_n_1121 = ~(mul_22_25_n_1079 | mul_22_25_n_1080);
 assign mul_22_25_n_1120 = ~(mul_22_25_n_1081 | mul_22_25_n_1082);
 assign mul_22_25_n_1119 = ~(mul_22_25_n_1079 & mul_22_25_n_1080);
 assign mul_22_25_n_1118 = ~(mul_22_25_n_1073 | mul_22_25_n_1076);
 assign mul_22_25_n_1117 = ~(mul_22_25_n_1077 & mul_22_25_n_1078);
 assign mul_22_25_n_1116 = ~(mul_22_25_n_1081 & mul_22_25_n_1082);
 assign mul_22_25_n_1115 = ~(mul_22_25_n_1071 | mul_22_25_n_1072);
 assign mul_22_25_n_1114 = ~(mul_22_25_n_1074 & mul_22_25_n_1075);
 assign mul_22_25_n_1113 = ~(mul_22_25_n_1071 & mul_22_25_n_1072);
 assign mul_22_25_n_1112 = ~(mul_22_25_n_1073 & mul_22_25_n_1076);
 assign mul_22_25_n_1111 = ~(mul_22_25_n_990 & mul_22_25_n_1053);
 assign mul_22_25_n_1110 = ~(mul_22_25_n_1083 & mul_22_25_n_1084);
 assign mul_22_25_n_1109 = ~(mul_22_25_n_1062 | mul_22_25_n_1085);
 assign mul_22_25_n_1108 = ~(mul_22_25_n_1069 & mul_22_25_n_1070);
 assign mul_22_25_n_1107 = ~(mul_22_25_n_1063 | mul_22_25_n_1064);
 assign mul_22_25_n_1106 = ~(mul_22_25_n_1077 | mul_22_25_n_1078);
 assign asc001_15_ = ~(mul_22_25_n_1031 ^ mul_22_25_n_1052);
 assign mul_22_25_n_1105 = ~(mul_22_25_n_1059 | n_119);
 assign mul_22_25_n_1104 = ~(mul_22_25_n_1774 & mul_22_25_n_1809);
 assign mul_22_25_n_1103 = ~(mul_22_25_n_1760 & mul_22_25_n_1795);
 assign mul_22_25_n_1102 = ~(mul_22_25_n_1057 | mul_22_25_n_1056);
 assign mul_22_25_n_1101 = ~(mul_22_25_n_1063 & mul_22_25_n_1064);
 assign mul_22_25_n_1100 = ~(mul_22_25_n_1761 & mul_22_25_n_1796);
 assign mul_22_25_n_1099 = ~(mul_22_25_n_1061 | n_51);
 assign mul_22_25_n_1098 = ~(mul_22_25_n_1058 | mul_22_25_n_1060);
 assign mul_22_25_n_1097 = ~(mul_22_25_n_1061 & n_51);
 assign mul_22_25_n_1096 = ~(mul_22_25_n_1065 & mul_22_25_n_1068);
 assign mul_22_25_n_1095 = ~(mul_22_25_n_1762 | mul_22_25_n_1797);
 assign mul_22_25_n_1094 = ~(mul_22_25_n_1059 & n_119);
 assign mul_22_25_n_1093 = ~(mul_22_25_n_1058 & mul_22_25_n_1060);
 assign mul_22_25_n_1092 = ~(mul_22_25_n_1761 | mul_22_25_n_1796);
 assign mul_22_25_n_1091 = ~(mul_22_25_n_1055 | mul_22_25_n_1054);
 assign mul_22_25_n_1090 = ~(mul_22_25_n_1057 & mul_22_25_n_1056);
 assign mul_22_25_n_1089 = ~(mul_22_25_n_990 | mul_22_25_n_1053);
 assign mul_22_25_n_1088 = ~(mul_22_25_n_1055 & mul_22_25_n_1054);
 assign mul_22_25_n_1087 = (mul_22_25_n_1062 & mul_22_25_n_1085);
 assign mul_22_25_n_1085 = ~mul_22_25_n_1798;
 assign mul_22_25_n_1084 = ~mul_22_25_n_1805;
 assign mul_22_25_n_1083 = ~mul_22_25_n_1770;
 assign mul_22_25_n_1082 = ~mul_22_25_n_1804;
 assign mul_22_25_n_1081 = ~mul_22_25_n_1769;
 assign mul_22_25_n_1080 = ~mul_22_25_n_1803;
 assign mul_22_25_n_1079 = ~mul_22_25_n_1768;
 assign mul_22_25_n_1078 = ~mul_22_25_n_1802;
 assign mul_22_25_n_1077 = ~mul_22_25_n_1767;
 assign mul_22_25_n_1076 = ~mul_22_25_n_1812;
 assign mul_22_25_n_1075 = ~mul_22_25_n_1801;
 assign mul_22_25_n_1074 = ~mul_22_25_n_1766;
 assign mul_22_25_n_1073 = ~mul_22_25_n_1777;
 assign mul_22_25_n_1072 = ~mul_22_25_n_1800;
 assign mul_22_25_n_1071 = ~mul_22_25_n_1765;
 assign mul_22_25_n_1070 = ~mul_22_25_n_1799;
 assign mul_22_25_n_1069 = ~mul_22_25_n_1764;
 assign mul_22_25_n_1068 = ~mul_22_25_n_1811;
 assign mul_22_25_n_1067 = ~(mul_22_25_n_1047 & (mul_22_25_n_1048 & (mul_22_25_n_980 | mul_22_25_n_1042)));
 assign mul_22_25_n_1066 = ~mul_22_25_n_1794;
 assign mul_22_25_n_1065 = ~mul_22_25_n_1776;
 assign mul_22_25_n_1064 = ~mul_22_25_n_1810;
 assign mul_22_25_n_1063 = ~mul_22_25_n_1775;
 assign mul_22_25_n_1062 = ~mul_22_25_n_1763;
 assign mul_22_25_n_1061 = ~mul_22_25_n_1759;
 assign mul_22_25_n_1060 = ~mul_22_25_n_1808;
 assign mul_22_25_n_1058 = ~mul_22_25_n_1773;
 assign mul_22_25_n_1057 = ~mul_22_25_n_1772;
 assign mul_22_25_n_1056 = ~mul_22_25_n_1807;
 assign mul_22_25_n_1055 = ~mul_22_25_n_1771;
 assign mul_22_25_n_1054 = ~mul_22_25_n_1806;
 assign mul_22_25_n_1053 = ~mul_22_25_n_1814;
 assign mul_22_25_n_1052 = ~(n_74 | (mul_22_25_n_1044 & n_75));
 assign asc001_14_ = ~(mul_22_25_n_1029 ^ mul_22_25_n_1044);
 assign mul_22_25_n_1050 = ~(~mul_22_25_n_1045 & mul_22_25_n_1046);
 assign mul_22_25_n_1049 = ~(mul_22_25_n_972 & (n_69 & (mul_22_25_n_1039 | mul_22_25_n_973)));
 assign mul_22_25_n_1048 = ~(mul_22_25_n_1025 | (n_92 | (mul_22_25_n_1038 & mul_22_25_n_1026)));
 assign mul_22_25_n_1047 = (mul_22_25_n_985 | mul_22_25_n_1042);
 assign mul_22_25_n_1046 = ~(n_120 & n_118);
 assign mul_22_25_n_1045 = ~(n_120 | n_118);
 assign mul_22_25_n_1044 = ~(~mul_22_25_n_1038 & (mul_22_25_n_988 | mul_22_25_n_1036));
 assign asc001_13_ = ~(mul_22_25_n_1030 ^ mul_22_25_n_999);
 assign mul_22_25_n_1042 = ~(~mul_22_25_n_1036 & mul_22_25_n_1026);
 assign mul_22_25_n_1041 = ~(mul_22_25_n_973 | mul_22_25_n_1035);
 assign mul_22_25_n_1040 = ~(n_116 & (n_109 | n_57));
 assign mul_22_25_n_1039 = ~(n_127 | (n_128 & n_114));
 assign mul_22_25_n_1038 = ~(n_77 & (n_76 | n_79));
 assign mul_22_25_n_1037 = ~mul_22_25_n_1793;
 assign mul_22_25_n_1034 = ~(n_108 & n_43);
 assign mul_22_25_n_1033 = ~(~n_109 & n_116);
 assign mul_22_25_n_1032 = ~(n_95 & n_57);
 assign mul_22_25_n_1031 = ~(n_93 | n_92);
 assign mul_22_25_n_1036 = (n_76 | n_78);
 assign mul_22_25_n_1030 = ~(n_76 | ~n_77);
 assign mul_22_25_n_1035 = ~(n_128 & n_115);
 assign mul_22_25_n_1029 = ~(n_75 & ~n_74);
 assign mul_22_25_n_1025 = ~(n_93 | ~n_74);
 assign mul_22_25_n_1024 = ~(n_115 & ~n_114);
 assign mul_22_25_n_1023 = ~(n_108 & n_110);
 assign mul_22_25_n_1022 = ~(~n_43 & n_68);
 assign mul_22_25_n_1021 = ~(n_61 & ~n_42);
 assign mul_22_25_n_1028 = ~(n_108 & n_68);
 assign mul_22_25_n_1027 = ~(n_109 | ~n_95);
 assign mul_22_25_n_1026 = ~(~n_75 | n_93);
 assign mul_22_25_n_1020 = ~(n_128 & ~n_127);
 assign mul_22_25_n_1019 = ~(mul_22_25_n_1782 & mul_22_25_n_1817);
 assign mul_22_25_n_1018 = ~(mul_22_25_n_1756 & mul_22_25_n_1791);
 assign mul_22_25_n_1017 = ~(mul_22_25_n_1752 | mul_22_25_n_1787);
 assign mul_22_25_n_1016 = ~(mul_22_25_n_998 & mul_22_25_n_997);
 assign mul_22_25_n_1015 = ~(mul_22_25_n_993 & mul_22_25_n_994);
 assign mul_22_25_n_1014 = ~(mul_22_25_n_989 | mul_22_25_n_995);
 assign mul_22_25_n_1013 = ~(mul_22_25_n_989 & mul_22_25_n_995);
 assign mul_22_25_n_1012 = ~(mul_22_25_n_998 | mul_22_25_n_997);
 assign mul_22_25_n_1011 = ~(mul_22_25_n_1755 & mul_22_25_n_1790);
 assign mul_22_25_n_1010 = ~(mul_22_25_n_957 & mul_22_25_n_996);
 assign asc001_11_ = (mul_22_25_n_975 ^ mul_22_25_n_987);
 assign asc001_12_ = ~(mul_22_25_n_986 ^ mul_22_25_n_988);
 assign mul_22_25_n_1009 = ~(mul_22_25_n_957 | mul_22_25_n_996);
 assign mul_22_25_n_999 = (n_79 & (mul_22_25_n_988 | n_78));
 assign mul_22_25_n_1008 = ~(mul_22_25_n_1752 & mul_22_25_n_1787);
 assign mul_22_25_n_1007 = ~(mul_22_25_n_993 | mul_22_25_n_994);
 assign mul_22_25_n_1006 = ~(mul_22_25_n_991 | mul_22_25_n_992);
 assign mul_22_25_n_1005 = ~(mul_22_25_n_1754 | mul_22_25_n_1789);
 assign mul_22_25_n_1004 = ~(mul_22_25_n_991 & mul_22_25_n_992);
 assign mul_22_25_n_1003 = (mul_22_25_n_1755 | mul_22_25_n_1790);
 assign mul_22_25_n_1002 = ~(mul_22_25_n_1756 | mul_22_25_n_1791);
 assign mul_22_25_n_998 = ~mul_22_25_n_1265;
 assign mul_22_25_n_997 = ~mul_22_25_n_1783;
 assign mul_22_25_n_996 = ~mul_22_25_n_1784;
 assign mul_22_25_n_995 = ~mul_22_25_n_1816;
 assign mul_22_25_n_994 = ~mul_22_25_n_1815;
 assign mul_22_25_n_993 = ~mul_22_25_n_1780;
 assign mul_22_25_n_992 = ~mul_22_25_n_1788;
 assign mul_22_25_n_991 = ~mul_22_25_n_1753;
 assign mul_22_25_n_990 = ~mul_22_25_n_1779;
 assign mul_22_25_n_989 = ~mul_22_25_n_1781;
 assign mul_22_25_n_988 = (mul_22_25_n_980 & mul_22_25_n_985);
 assign mul_22_25_n_987 = ~(n_131 & (mul_22_25_n_982 | n_72));
 assign mul_22_25_n_986 = ~(~n_79 | n_78);
 assign mul_22_25_n_985 = ~(mul_22_25_n_976 | (n_71 | (n_63 & mul_22_25_n_978)));
 assign mul_22_25_n_984 = ~(mul_22_25_n_1751 & mul_22_25_n_1271);
 assign mul_22_25_n_983 = ~(mul_22_25_n_1751 | mul_22_25_n_1271);
 assign mul_22_25_n_982 = ~(n_146 | n_63);
 assign asc001_9_ = ~(n_62 ^ n_145);
 assign mul_22_25_n_980 = ~(n_146 & mul_22_25_n_978);
 assign mul_22_25_n_979 = ~(mul_22_25_n_967 & (mul_22_25_n_966 | mul_22_25_n_947));
 assign mul_22_25_n_976 = ~(n_44 | n_131);
 assign mul_22_25_n_978 = ~(n_44 | n_72);
 assign mul_22_25_n_977 = ~(mul_22_25_n_951 | mul_22_25_n_966);
 assign mul_22_25_n_975 = ~(n_44 | n_71);
 assign mul_22_25_n_974 = ~(n_72 | ~n_131);
 assign mul_22_25_n_972 = ~(n_45 & n_102);
 assign mul_22_25_n_971 = ~(mul_22_25_n_966 | ~mul_22_25_n_967);
 assign mul_22_25_n_970 = ~(n_138 & ~n_139);
 assign mul_22_25_n_969 = ~(n_45 & n_69);
 assign mul_22_25_n_968 = ~(~n_102 & n_103);
 assign mul_22_25_n_973 = ~(n_45 & n_103);
 assign mul_22_25_n_967 = ~(mul_22_25_n_1748 & mul_22_25_n_1786);
 assign mul_22_25_n_966 = ~(mul_22_25_n_1748 | mul_22_25_n_1786);
 assign mul_22_25_n_965 = ~(mul_22_25_n_1750 | mul_22_25_n_1272);
 assign mul_22_25_n_964 = ~(mul_22_25_n_1749 | mul_22_25_n_1273);
 assign mul_22_25_n_963 = ~(mul_22_25_n_1749 & mul_22_25_n_1273);
 assign mul_22_25_n_962 = ~(mul_22_25_n_933 | mul_22_25_n_952);
 assign mul_22_25_n_961 = ~(mul_22_25_n_1266 & mul_22_25_n_1269);
 assign mul_22_25_n_960 = ~(mul_22_25_n_933 & mul_22_25_n_952);
 assign mul_22_25_n_959 = ~(mul_22_25_n_954 & mul_22_25_n_953);
 assign mul_22_25_n_958 = ~(mul_22_25_n_954 | mul_22_25_n_953);
 assign mul_22_25_n_957 = ~mul_22_25_n_1818;
 assign asc001_8_ = ~(mul_22_25_n_950 ^ mul_22_25_n_949);
 assign mul_22_25_n_955 = (mul_22_25_n_951 & mul_22_25_n_947);
 assign mul_22_25_n_954 = ~mul_22_25_n_1268;
 assign mul_22_25_n_953 = ~mul_22_25_n_1270;
 assign mul_22_25_n_952 = ~mul_22_25_n_1267;
 assign mul_22_25_n_951 = ~(~mul_22_25_n_949 & mul_22_25_n_946);
 assign mul_22_25_n_950 = (mul_22_25_n_946 & mul_22_25_n_947);
 assign mul_22_25_n_949 = ~(mul_22_25_n_943 | (mul_22_25_n_944 | (mul_22_25_n_930 & mul_22_25_n_941)));
 assign asc001_7_ = (mul_22_25_n_940 ^ mul_22_25_n_942);
 assign mul_22_25_n_947 = ~(mul_22_25_n_1276 & mul_22_25_n_1278);
 assign mul_22_25_n_946 = (mul_22_25_n_1276 | mul_22_25_n_1278);
 assign asc001_6_ = ~(mul_22_25_n_932 ^ mul_22_25_n_939);
 assign mul_22_25_n_944 = (mul_22_25_n_929 & mul_22_25_n_941);
 assign mul_22_25_n_943 = ~(mul_22_25_n_937 & (mul_22_25_n_935 | mul_22_25_n_936));
 assign mul_22_25_n_942 = ~(mul_22_25_n_936 & (mul_22_25_n_932 | mul_22_25_n_934));
 assign mul_22_25_n_941 = ~(mul_22_25_n_935 | mul_22_25_n_934);
 assign mul_22_25_n_940 = ~(~mul_22_25_n_937 | mul_22_25_n_935);
 assign mul_22_25_n_939 = ~(mul_22_25_n_934 | ~mul_22_25_n_936);
 assign mul_22_25_n_938 = ~(mul_22_25_n_1274 ^ mul_22_25_n_1275);
 assign mul_22_25_n_937 = ~(mul_22_25_n_1277 & mul_22_25_n_1280);
 assign mul_22_25_n_936 = ~(mul_22_25_n_1279 & mul_22_25_n_1785);
 assign mul_22_25_n_935 = ~(mul_22_25_n_1277 | mul_22_25_n_1280);
 assign mul_22_25_n_934 = ~(mul_22_25_n_1279 | mul_22_25_n_1785);
 assign mul_22_25_n_933 = ~mul_22_25_n_1819;
 assign asc001_5_ = ~(mul_22_25_n_924 ^ mul_22_25_n_928);
 assign mul_22_25_n_932 = ~(mul_22_25_n_929 | mul_22_25_n_930);
 assign mul_22_25_n_930 = ~(mul_22_25_n_927 & (mul_22_25_n_921 | mul_22_25_n_926));
 assign mul_22_25_n_929 = ~(mul_22_25_n_922 | mul_22_25_n_926);
 assign mul_22_25_n_928 = ~(mul_22_25_n_926 | ~mul_22_25_n_927);
 assign mul_22_25_n_927 = ~(mul_22_25_n_1281 & mul_22_25_n_1283);
 assign mul_22_25_n_926 = ~(mul_22_25_n_1281 | mul_22_25_n_1283);
 assign asc001_4_ = ~(mul_22_25_n_919 ^ mul_22_25_n_923);
 assign mul_22_25_n_924 = (mul_22_25_n_922 & mul_22_25_n_921);
 assign mul_22_25_n_923 = ~(mul_22_25_n_921 & mul_22_25_n_920);
 assign mul_22_25_n_922 = ~(mul_22_25_n_919 & mul_22_25_n_920);
 assign mul_22_25_n_921 = ~(mul_22_25_n_889 & mul_22_25_n_1282);
 assign mul_22_25_n_920 = (mul_22_25_n_889 | mul_22_25_n_1282);
 assign asc001_3_ = ~(mul_22_25_n_915 ^ mul_22_25_n_916);
 assign mul_22_25_n_919 = ~(mul_22_25_n_917 & (mul_22_25_n_913 & (mul_22_25_n_914 | mul_22_25_n_911)));
 assign mul_22_25_n_917 = ~(mul_22_25_n_833 & ~mul_22_25_n_914);
 assign mul_22_25_n_916 = ~(mul_22_25_n_913 & ~mul_22_25_n_914);
 assign mul_22_25_n_915 = ~(~mul_22_25_n_833 & mul_22_25_n_911);
 assign mul_22_25_n_914 = ~(mul_22_25_n_900 | mul_22_25_n_849);
 assign mul_22_25_n_913 = ~(mul_22_25_n_900 & mul_22_25_n_849);
 assign asc001_2_ = ~(mul_22_25_n_830 ^ mul_22_25_n_879);
 assign mul_22_25_n_911 = ~(mul_22_25_n_864 & mul_22_25_n_830);
 assign mul_22_25_n_910 = ~(mul_22_25_n_878 & (mul_22_25_n_858 | mul_22_25_n_711));
 assign mul_22_25_n_909 = (mul_22_25_n_847 ^ mul_22_25_n_535);
 assign mul_22_25_n_908 = (mul_22_25_n_533 ^ mul_22_25_n_845);
 assign mul_22_25_n_907 = (mul_22_25_n_538 ^ mul_22_25_n_832);
 assign mul_22_25_n_906 = ~(mul_22_25_n_559 ^ mul_22_25_n_831);
 assign mul_22_25_n_905 = ~(mul_22_25_n_836 ^ mul_22_25_n_839);
 assign mul_22_25_n_904 = (n_210 ^ mul_22_25_n_846);
 assign mul_22_25_n_903 = ~(mul_22_25_n_560 ^ mul_22_25_n_707);
 assign mul_22_25_n_902 = (mul_22_25_n_558 ^ mul_22_25_n_705);
 assign mul_22_25_n_901 = (mul_22_25_n_556 ^ mul_22_25_n_844);
 assign mul_22_25_n_899 = (mul_22_25_n_835 ^ mul_22_25_n_557);
 assign mul_22_25_n_898 = (mul_22_25_n_536 ^ mul_22_25_n_710);
 assign mul_22_25_n_897 = ~(mul_22_25_n_534 ^ mul_22_25_n_706);
 assign mul_22_25_n_896 = (mul_22_25_n_838 ^ mul_22_25_n_709);
 assign mul_22_25_n_895 = (mul_22_25_n_834 ^ mul_22_25_n_531);
 assign mul_22_25_n_894 = (mul_22_25_n_539 ^ mul_22_25_n_708);
 assign mul_22_25_n_893 = (mul_22_25_n_532 ^ mul_22_25_n_848);
 assign mul_22_25_n_892 = (mul_22_25_n_540 ^ mul_22_25_n_842);
 assign mul_22_25_n_891 = (mul_22_25_n_840 ^ mul_22_25_n_541);
 assign mul_22_25_n_890 = (mul_22_25_n_841 ^ mul_22_25_n_555);
 assign mul_22_25_n_900 = (mul_22_25_n_537 ^ mul_22_25_n_837);
 assign mul_22_25_n_888 = ~(mul_22_25_n_541 | mul_22_25_n_840);
 assign mul_22_25_n_887 = ~(mul_22_25_n_540 | mul_22_25_n_842);
 assign mul_22_25_n_886 = ~(mul_22_25_n_557 | mul_22_25_n_835);
 assign mul_22_25_n_885 = ~(mul_22_25_n_532 | mul_22_25_n_848);
 assign mul_22_25_n_884 = ~(mul_22_25_n_709 | mul_22_25_n_838);
 assign mul_22_25_n_883 = ~(mul_22_25_n_531 | mul_22_25_n_834);
 assign mul_22_25_n_882 = ~(mul_22_25_n_555 | mul_22_25_n_841);
 assign mul_22_25_n_881 = ~(mul_22_25_n_836 | ~mul_22_25_n_839);
 assign mul_22_25_n_880 = ~(mul_22_25_n_846 | n_210);
 assign mul_22_25_n_879 = ~(mul_22_25_n_864 & ~mul_22_25_n_833);
 assign mul_22_25_n_889 = ~(mul_22_25_n_537 | mul_22_25_n_837);
 assign mul_22_25_n_877 = ~(mul_22_25_n_560 | ~mul_22_25_n_707);
 assign mul_22_25_n_876 = ~(mul_22_25_n_847 | mul_22_25_n_535);
 assign mul_22_25_n_875 = ~(mul_22_25_n_845 | mul_22_25_n_533);
 assign mul_22_25_n_874 = ~(mul_22_25_n_832 | mul_22_25_n_538);
 assign mul_22_25_n_873 = ~(mul_22_25_n_710 | mul_22_25_n_536);
 assign mul_22_25_n_872 = ~(mul_22_25_n_708 | mul_22_25_n_539);
 assign mul_22_25_n_871 = ~(mul_22_25_n_534 | ~mul_22_25_n_706);
 assign mul_22_25_n_870 = ~(mul_22_25_n_705 | mul_22_25_n_558);
 assign mul_22_25_n_869 = ~(mul_22_25_n_844 | mul_22_25_n_556);
 assign mul_22_25_n_868 = ~(mul_22_25_n_831 | ~mul_22_25_n_559);
 assign asc001_1_ = ~(mul_22_25_n_830 | (mul_22_25_n_561 & mul_22_25_n_447));
 assign mul_22_25_n_878 = ~(mul_22_25_n_858 & mul_22_25_n_711);
 assign mul_22_25_n_866 = ~mul_22_25_n_865;
 assign mul_22_25_n_863 = ~mul_22_25_n_862;
 assign mul_22_25_n_861 = ~mul_22_25_n_860;
 assign mul_22_25_n_859 = ~mul_22_25_n_0;
 assign mul_22_25_n_857 = ~mul_22_25_n_856;
 assign mul_22_25_n_855 = ~mul_22_25_n_854;
 assign mul_22_25_n_853 = ~mul_22_25_n_852;
 assign mul_22_25_n_851 = ~mul_22_25_n_850;
 assign mul_22_25_n_829 = ~((mul_22_25_n_280 | mul_22_25_n_221) & (mul_22_25_n_485 | mul_22_25_n_376));
 assign mul_22_25_n_828 = ~((mul_22_25_n_281 | mul_22_25_n_253) & (mul_22_25_n_493 | mul_22_25_n_390));
 assign mul_22_25_n_827 = ~((mul_22_25_n_284 | mul_22_25_n_403) & (mul_22_25_n_491 | mul_22_25_n_442));
 assign mul_22_25_n_826 = ~((mul_22_25_n_285 | mul_22_25_n_364) & (mul_22_25_n_489 | mul_22_25_n_314));
 assign mul_22_25_n_825 = ~((mul_22_25_n_286 | mul_22_25_n_290) & (mul_22_25_n_483 | mul_22_25_n_242));
 assign mul_22_25_n_824 = ~((mul_22_25_n_287 | mul_22_25_n_362) & (mul_22_25_n_479 | mul_22_25_n_402));
 assign mul_22_25_n_823 = ~((mul_22_25_n_280 | mul_22_25_n_368) & (mul_22_25_n_485 | mul_22_25_n_135));
 assign mul_22_25_n_822 = ~((mul_22_25_n_282 | mul_22_25_n_111) & (mul_22_25_n_481 | mul_22_25_n_216));
 assign mul_22_25_n_821 = ~((mul_22_25_n_284 | mul_22_25_n_106) & (mul_22_25_n_491 | mul_22_25_n_254));
 assign mul_22_25_n_820 = ~((mul_22_25_n_283 | mul_22_25_n_126) & (mul_22_25_n_487 | mul_22_25_n_164));
 assign mul_22_25_n_819 = ~((mul_22_25_n_280 | mul_22_25_n_217) & (mul_22_25_n_485 | mul_22_25_n_227));
 assign mul_22_25_n_818 = ~((mul_22_25_n_280 | mul_22_25_n_376) & (mul_22_25_n_485 | mul_22_25_n_267));
 assign mul_22_25_n_817 = ~((mul_22_25_n_283 | mul_22_25_n_411) & (mul_22_25_n_487 | mul_22_25_n_344));
 assign mul_22_25_n_816 = ~((mul_22_25_n_287 | mul_22_25_n_246) & (mul_22_25_n_479 | mul_22_25_n_244));
 assign mul_22_25_n_815 = ~(mul_22_25_n_519 | (mul_22_25_n_486 & mul_22_25_n_418));
 assign mul_22_25_n_814 = ~((mul_22_25_n_283 | mul_22_25_n_366) & (mul_22_25_n_487 | mul_22_25_n_371));
 assign mul_22_25_n_813 = ~(mul_22_25_n_520 | (mul_22_25_n_490 & mul_22_25_n_438));
 assign mul_22_25_n_812 = ~((mul_22_25_n_285 | mul_22_25_n_143) & (mul_22_25_n_489 | mul_22_25_n_324));
 assign mul_22_25_n_811 = ~(mul_22_25_n_3 | (mul_22_25_n_488 & mul_22_25_n_429));
 assign mul_22_25_n_810 = ~(mul_22_25_n_521 & (mul_22_25_n_485 | mul_22_25_n_437));
 assign mul_22_25_n_809 = ~(mul_22_25_n_515 | (mul_22_25_n_480 & mul_22_25_n_420));
 assign mul_22_25_n_808 = ~(mul_22_25_n_2 & (mul_22_25_n_487 | mul_22_25_n_434));
 assign mul_22_25_n_807 = ~(mul_22_25_n_5 | (mul_22_25_n_482 & mul_22_25_n_417));
 assign mul_22_25_n_806 = ~((mul_22_25_n_286 | mul_22_25_n_265) & (mul_22_25_n_483 | mul_22_25_n_226));
 assign mul_22_25_n_805 = ~(mul_22_25_n_518 | (mul_22_25_n_478 & mul_22_25_n_431));
 assign mul_22_25_n_804 = ~((mul_22_25_n_287 | mul_22_25_n_255) & (mul_22_25_n_479 | mul_22_25_n_338));
 assign mul_22_25_n_803 = ~((mul_22_25_n_288 | mul_22_25_n_270) & (mul_22_25_n_494 | mul_22_25_n_436));
 assign mul_22_25_n_802 = ~((mul_22_25_n_280 | mul_22_25_n_407) & (mul_22_25_n_485 | mul_22_25_n_100));
 assign mul_22_25_n_801 = ~((mul_22_25_n_282 | mul_22_25_n_198) & (mul_22_25_n_481 | mul_22_25_n_98));
 assign mul_22_25_n_800 = ~((mul_22_25_n_283 | mul_22_25_n_164) & (mul_22_25_n_487 | mul_22_25_n_103));
 assign mul_22_25_n_799 = ~((mul_22_25_n_288 | mul_22_25_n_155) & (mul_22_25_n_494 | mul_22_25_n_96));
 assign mul_22_25_n_798 = ~((mul_22_25_n_285 | mul_22_25_n_292) & (mul_22_25_n_489 | mul_22_25_n_104));
 assign mul_22_25_n_797 = ~((mul_22_25_n_284 | mul_22_25_n_291) & (mul_22_25_n_491 | mul_22_25_n_97));
 assign mul_22_25_n_796 = ~((mul_22_25_n_288 | mul_22_25_n_404) & (mul_22_25_n_494 | mul_22_25_n_155));
 assign mul_22_25_n_795 = ~((mul_22_25_n_287 | mul_22_25_n_241) & (mul_22_25_n_479 | mul_22_25_n_101));
 assign mul_22_25_n_794 = ~((mul_22_25_n_286 | mul_22_25_n_317) & (mul_22_25_n_483 | mul_22_25_n_95));
 assign mul_22_25_n_793 = ~((mul_22_25_n_282 | mul_22_25_n_330) & (mul_22_25_n_481 | mul_22_25_n_180));
 assign mul_22_25_n_792 = ~((mul_22_25_n_286 | mul_22_25_n_414) & (mul_22_25_n_483 | mul_22_25_n_384));
 assign mul_22_25_n_791 = ~((mul_22_25_n_286 | mul_22_25_n_308) & (mul_22_25_n_483 | mul_22_25_n_410));
 assign mul_22_25_n_790 = ~((mul_22_25_n_287 | mul_22_25_n_124) & (mul_22_25_n_479 | mul_22_25_n_122));
 assign mul_22_25_n_789 = ~((mul_22_25_n_284 | mul_22_25_n_333) & (mul_22_25_n_491 | mul_22_25_n_186));
 assign mul_22_25_n_788 = ~((mul_22_25_n_288 | mul_22_25_n_163) & (mul_22_25_n_494 | mul_22_25_n_295));
 assign mul_22_25_n_787 = ~((mul_22_25_n_286 | mul_22_25_n_242) & (mul_22_25_n_483 | mul_22_25_n_207));
 assign mul_22_25_n_786 = ~((mul_22_25_n_288 | mul_22_25_n_158) & (mul_22_25_n_494 | mul_22_25_n_369));
 assign mul_22_25_n_785 = ~((mul_22_25_n_288 | mul_22_25_n_266) & (mul_22_25_n_494 | mul_22_25_n_131));
 assign mul_22_25_n_784 = ~((mul_22_25_n_283 | mul_22_25_n_231) & (mul_22_25_n_487 | mul_22_25_n_181));
 assign mul_22_25_n_783 = ~((mul_22_25_n_285 | mul_22_25_n_252) & (mul_22_25_n_489 | mul_22_25_n_336));
 assign mul_22_25_n_782 = ~((mul_22_25_n_283 | mul_22_25_n_148) & (mul_22_25_n_487 | mul_22_25_n_378));
 assign mul_22_25_n_781 = ~((mul_22_25_n_280 | mul_22_25_n_379) & (mul_22_25_n_485 | mul_22_25_n_249));
 assign mul_22_25_n_780 = ~((mul_22_25_n_285 | mul_22_25_n_225) & (mul_22_25_n_489 | mul_22_25_n_145));
 assign mul_22_25_n_779 = ~((mul_22_25_n_281 | mul_22_25_n_175) & (mul_22_25_n_493 | mul_22_25_n_237));
 assign mul_22_25_n_778 = ~((mul_22_25_n_280 | mul_22_25_n_141) & (mul_22_25_n_485 | mul_22_25_n_413));
 assign mul_22_25_n_777 = ~((mul_22_25_n_281 | mul_22_25_n_387) & (mul_22_25_n_493 | mul_22_25_n_406));
 assign mul_22_25_n_776 = ~((mul_22_25_n_287 | mul_22_25_n_347) & (mul_22_25_n_479 | mul_22_25_n_189));
 assign mul_22_25_n_775 = ~((mul_22_25_n_284 | mul_22_25_n_173) & (mul_22_25_n_491 | mul_22_25_n_139));
 assign mul_22_25_n_774 = ~((mul_22_25_n_284 | mul_22_25_n_395) & (mul_22_25_n_491 | mul_22_25_n_391));
 assign mul_22_25_n_773 = ~((mul_22_25_n_286 | mul_22_25_n_433) & (mul_22_25_n_483 | mul_22_25_n_372));
 assign mul_22_25_n_772 = ~((mul_22_25_n_282 | mul_22_25_n_337) & (mul_22_25_n_481 | mul_22_25_n_409));
 assign mul_22_25_n_771 = ~((mul_22_25_n_285 | mul_22_25_n_314) & (mul_22_25_n_489 | mul_22_25_n_215));
 assign mul_22_25_n_770 = ~((mul_22_25_n_284 | mul_22_25_n_318) & (mul_22_25_n_491 | mul_22_25_n_415));
 assign mul_22_25_n_769 = ~((mul_22_25_n_286 | mul_22_25_n_329) & (mul_22_25_n_483 | mul_22_25_n_317));
 assign mul_22_25_n_768 = ~((mul_22_25_n_287 | mul_22_25_n_359) & (mul_22_25_n_479 | mul_22_25_n_241));
 assign mul_22_25_n_767 = ~((mul_22_25_n_288 | mul_22_25_n_121) & (mul_22_25_n_494 | mul_22_25_n_177));
 assign mul_22_25_n_766 = ~((mul_22_25_n_283 | mul_22_25_n_394) & (mul_22_25_n_487 | mul_22_25_n_148));
 assign mul_22_25_n_765 = ~((mul_22_25_n_285 | mul_22_25_n_419) & (mul_22_25_n_489 | mul_22_25_n_127));
 assign mul_22_25_n_764 = ~((mul_22_25_n_280 | mul_22_25_n_296) & (mul_22_25_n_485 | mul_22_25_n_379));
 assign mul_22_25_n_763 = ~((mul_22_25_n_280 | mul_22_25_n_437) & (mul_22_25_n_485 | mul_22_25_n_248));
 assign mul_22_25_n_762 = ~((mul_22_25_n_285 | mul_22_25_n_399) & (mul_22_25_n_489 | mul_22_25_n_219));
 assign mul_22_25_n_761 = ~((mul_22_25_n_281 | mul_22_25_n_390) & (mul_22_25_n_493 | mul_22_25_n_299));
 assign mul_22_25_n_760 = ~((mul_22_25_n_280 | mul_22_25_n_133) & (mul_22_25_n_485 | mul_22_25_n_298));
 assign mul_22_25_n_759 = ~((mul_22_25_n_285 | mul_22_25_n_373) & (mul_22_25_n_489 | mul_22_25_n_252));
 assign mul_22_25_n_758 = ~((mul_22_25_n_283 | mul_22_25_n_441) & (mul_22_25_n_487 | mul_22_25_n_190));
 assign mul_22_25_n_757 = ~((mul_22_25_n_280 | mul_22_25_n_413) & (mul_22_25_n_485 | mul_22_25_n_263));
 assign mul_22_25_n_756 = ~((mul_22_25_n_287 | mul_22_25_n_352) & (mul_22_25_n_479 | mul_22_25_n_184));
 assign mul_22_25_n_755 = ~((mul_22_25_n_287 | mul_22_25_n_402) & (mul_22_25_n_479 | mul_22_25_n_110));
 assign mul_22_25_n_754 = ~((mul_22_25_n_285 | mul_22_25_n_423) & (mul_22_25_n_489 | mul_22_25_n_143));
 assign mul_22_25_n_753 = ~((mul_22_25_n_286 | mul_22_25_n_136) & (mul_22_25_n_483 | mul_22_25_n_375));
 assign mul_22_25_n_752 = ~((mul_22_25_n_286 | mul_22_25_n_226) & (mul_22_25_n_483 | mul_22_25_n_446));
 assign mul_22_25_n_751 = ~((mul_22_25_n_282 | mul_22_25_n_448) & (mul_22_25_n_481 | mul_22_25_n_377));
 assign mul_22_25_n_750 = ~((mul_22_25_n_286 | mul_22_25_n_382) & (mul_22_25_n_483 | mul_22_25_n_196));
 assign mul_22_25_n_749 = ~((mul_22_25_n_287 | mul_22_25_n_238) & (mul_22_25_n_479 | mul_22_25_n_354));
 assign mul_22_25_n_748 = ~((mul_22_25_n_288 | mul_22_25_n_370) & (mul_22_25_n_494 | mul_22_25_n_348));
 assign mul_22_25_n_747 = ~((mul_22_25_n_281 | mul_22_25_n_445) & (mul_22_25_n_493 | mul_22_25_n_257));
 assign mul_22_25_n_746 = ~((mul_22_25_n_285 | mul_22_25_n_130) & (mul_22_25_n_489 | mul_22_25_n_373));
 assign mul_22_25_n_745 = ~((mul_22_25_n_283 | mul_22_25_n_360) & (mul_22_25_n_487 | mul_22_25_n_394));
 assign mul_22_25_n_744 = ~((mul_22_25_n_280 | mul_22_25_n_135) & (mul_22_25_n_485 | mul_22_25_n_296));
 assign mul_22_25_n_743 = ~((mul_22_25_n_287 | mul_22_25_n_189) & (mul_22_25_n_479 | mul_22_25_n_255));
 assign mul_22_25_n_742 = ~((mul_22_25_n_282 | mul_22_25_n_168) & (mul_22_25_n_481 | mul_22_25_n_325));
 assign mul_22_25_n_741 = ~((mul_22_25_n_282 | mul_22_25_n_156) & (mul_22_25_n_481 | mul_22_25_n_313));
 assign mul_22_25_n_740 = ~((mul_22_25_n_288 | mul_22_25_n_348) & (mul_22_25_n_494 | mul_22_25_n_266));
 assign mul_22_25_n_739 = ~((mul_22_25_n_284 | mul_22_25_n_139) & (mul_22_25_n_491 | mul_22_25_n_106));
 assign mul_22_25_n_738 = ~((mul_22_25_n_283 | mul_22_25_n_381) & (mul_22_25_n_487 | mul_22_25_n_366));
 assign mul_22_25_n_737 = ~((mul_22_25_n_283 | mul_22_25_n_233) & (mul_22_25_n_487 | mul_22_25_n_126));
 assign mul_22_25_n_736 = ~((mul_22_25_n_286 | mul_22_25_n_410) & (mul_22_25_n_483 | mul_22_25_n_112));
 assign mul_22_25_n_735 = ~((mul_22_25_n_285 | mul_22_25_n_332) & (mul_22_25_n_489 | mul_22_25_n_230));
 assign mul_22_25_n_734 = ~((mul_22_25_n_287 | mul_22_25_n_354) & (mul_22_25_n_479 | mul_22_25_n_124));
 assign mul_22_25_n_733 = ~((mul_22_25_n_287 | mul_22_25_n_338) & (mul_22_25_n_479 | mul_22_25_n_352));
 assign mul_22_25_n_732 = ~((mul_22_25_n_287 | mul_22_25_n_235) & (mul_22_25_n_479 | mul_22_25_n_238));
 assign mul_22_25_n_731 = ~((mul_22_25_n_288 | mul_22_25_n_392) & (mul_22_25_n_494 | mul_22_25_n_370));
 assign mul_22_25_n_730 = ~((mul_22_25_n_283 | mul_22_25_n_344) & (mul_22_25_n_487 | mul_22_25_n_231));
 assign mul_22_25_n_729 = ~((mul_22_25_n_285 | mul_22_25_n_223) & (mul_22_25_n_489 | mul_22_25_n_130));
 assign mul_22_25_n_728 = ~((mul_22_25_n_285 | mul_22_25_n_250) & (mul_22_25_n_489 | mul_22_25_n_399));
 assign mul_22_25_n_727 = ~((mul_22_25_n_284 | mul_22_25_n_254) & (mul_22_25_n_491 | mul_22_25_n_182));
 assign mul_22_25_n_726 = ~((mul_22_25_n_282 | mul_22_25_n_313) & (mul_22_25_n_481 | mul_22_25_n_337));
 assign mul_22_25_n_725 = ~((mul_22_25_n_284 | mul_22_25_n_335) & (mul_22_25_n_491 | mul_22_25_n_318));
 assign mul_22_25_n_724 = ~((mul_22_25_n_285 | mul_22_25_n_302) & (mul_22_25_n_489 | mul_22_25_n_250));
 assign mul_22_25_n_723 = ~((mul_22_25_n_284 | mul_22_25_n_259) & (mul_22_25_n_491 | mul_22_25_n_335));
 assign mul_22_25_n_722 = ~((mul_22_25_n_281 | mul_22_25_n_264) & (mul_22_25_n_493 | mul_22_25_n_256));
 assign mul_22_25_n_721 = ~((mul_22_25_n_280 | mul_22_25_n_267) & (mul_22_25_n_485 | mul_22_25_n_368));
 assign mul_22_25_n_720 = ~((mul_22_25_n_284 | mul_22_25_n_311) & (mul_22_25_n_491 | mul_22_25_n_331));
 assign mul_22_25_n_719 = ~((mul_22_25_n_286 | mul_22_25_n_446) & (mul_22_25_n_483 | mul_22_25_n_414));
 assign mul_22_25_n_718 = ~((mul_22_25_n_287 | mul_22_25_n_303) & (mul_22_25_n_479 | mul_22_25_n_416));
 assign mul_22_25_n_717 = ~((mul_22_25_n_282 | mul_22_25_n_444) & (mul_22_25_n_481 | mul_22_25_n_304));
 assign mul_22_25_n_716 = ~((mul_22_25_n_286 | mul_22_25_n_207) & (mul_22_25_n_483 | mul_22_25_n_265));
 assign mul_22_25_n_715 = ~((mul_22_25_n_283 | mul_22_25_n_193) & (mul_22_25_n_487 | mul_22_25_n_159));
 assign mul_22_25_n_714 = ~((mul_22_25_n_281 | mul_22_25_n_165) & (mul_22_25_n_493 | mul_22_25_n_120));
 assign mul_22_25_n_713 = ~((mul_22_25_n_285 | mul_22_25_n_324) & (mul_22_25_n_489 | mul_22_25_n_223));
 assign mul_22_25_n_712 = ~((mul_22_25_n_283 | mul_22_25_n_371) & (mul_22_25_n_487 | mul_22_25_n_218));
 assign mul_22_25_n_865 = ~(mul_22_25_n_517 & (mul_22_25_n_493 | mul_22_25_n_425));
 assign mul_22_25_n_864 = ~(mul_22_25_n_542 & mul_22_25_n_516);
 assign mul_22_25_n_862 = ~((mul_22_25_n_457 & mul_22_25_n_247) | (mul_22_25_n_484 & mul_22_25_n_356));
 assign mul_22_25_n_860 = ~(mul_22_25_n_4 & (mul_22_25_n_479 | mul_22_25_n_422));
 assign mul_22_25_n_858 = ~((mul_22_25_n_455 & mul_22_25_n_426) | (mul_22_25_n_492 & mul_22_25_n_341));
 assign mul_22_25_n_856 = ~((mul_22_25_n_454 & mul_22_25_n_289) | (mul_22_25_n_480 & mul_22_25_n_229));
 assign mul_22_25_n_854 = ~(mul_22_25_n_515 | (mul_22_25_n_480 & mul_22_25_n_427));
 assign mul_22_25_n_852 = ~(mul_22_25_n_5 | (mul_22_25_n_482 & mul_22_25_n_432));
 assign mul_22_25_n_850 = ~(mul_22_25_n_520 | (mul_22_25_n_490 & mul_22_25_n_428));
 assign mul_22_25_n_849 = ~((mul_22_25_n_281 | mul_22_25_n_214) & (mul_22_25_n_493 | mul_22_25_n_102));
 assign mul_22_25_n_848 = ~(mul_22_25_n_545 & {in1[5]});
 assign mul_22_25_n_847 = ~((mul_22_25_n_455 & mul_22_25_n_211) | (mul_22_25_n_492 & mul_22_25_n_154));
 assign mul_22_25_n_846 = ~((mul_22_25_n_455 & mul_22_25_n_305) | (mul_22_25_n_492 & mul_22_25_n_174));
 assign mul_22_25_n_845 = ~((mul_22_25_n_455 & mul_22_25_n_144) | (mul_22_25_n_492 & mul_22_25_n_211));
 assign mul_22_25_n_844 = ~((mul_22_25_n_455 & mul_22_25_n_161) | (mul_22_25_n_492 & mul_22_25_n_385));
 assign mul_22_25_n_842 = ~(mul_22_25_n_546 & {in1[17]});
 assign mul_22_25_n_841 = ~(mul_22_25_n_548 & {in1[15]});
 assign mul_22_25_n_840 = ~(mul_22_25_n_549 & {in1[7]});
 assign mul_22_25_n_839 = ~((mul_22_25_n_281 | mul_22_25_n_257) & (mul_22_25_n_493 | mul_22_25_n_387));
 assign mul_22_25_n_838 = ~(mul_22_25_n_551 & {in1[9]});
 assign mul_22_25_n_837 = ~(mul_22_25_n_552 & {in1[3]});
 assign mul_22_25_n_836 = ~(mul_22_25_n_550 & {in1[11]});
 assign mul_22_25_n_835 = ~(mul_22_25_n_553 & {in1[19]});
 assign mul_22_25_n_834 = ~(mul_22_25_n_547 & {in1[13]});
 assign mul_22_25_n_833 = ~(mul_22_25_n_542 | mul_22_25_n_516);
 assign mul_22_25_n_832 = ~((mul_22_25_n_455 & mul_22_25_n_232) | (mul_22_25_n_492 & mul_22_25_n_144));
 assign mul_22_25_n_831 = ~((mul_22_25_n_455 & mul_22_25_n_341) | (mul_22_25_n_492 & mul_22_25_n_232));
 assign mul_22_25_n_830 = ~(mul_22_25_n_561 | mul_22_25_n_447);
 assign mul_22_25_n_704 = ~((mul_22_25_n_288 | mul_22_25_n_295) & (mul_22_25_n_494 | mul_22_25_n_392));
 assign mul_22_25_n_703 = ~((mul_22_25_n_287 | mul_22_25_n_309) & (mul_22_25_n_479 | mul_22_25_n_246));
 assign mul_22_25_n_702 = ~((mul_22_25_n_286 | mul_22_25_n_258) & (mul_22_25_n_483 | mul_22_25_n_308));
 assign mul_22_25_n_701 = ~((mul_22_25_n_282 | mul_22_25_n_114) & (mul_22_25_n_481 | mul_22_25_n_116));
 assign mul_22_25_n_700 = ~((mul_22_25_n_286 | mul_22_25_n_204) & (mul_22_25_n_483 | mul_22_25_n_382));
 assign mul_22_25_n_699 = ~((mul_22_25_n_288 | mul_22_25_n_326) & (mul_22_25_n_494 | mul_22_25_n_199));
 assign mul_22_25_n_698 = ~((mul_22_25_n_281 | mul_22_25_n_299) & (mul_22_25_n_493 | mul_22_25_n_445));
 assign mul_22_25_n_697 = ~((mul_22_25_n_288 | mul_22_25_n_203) & (mul_22_25_n_494 | mul_22_25_n_151));
 assign mul_22_25_n_696 = ~((mul_22_25_n_285 | mul_22_25_n_215) & (mul_22_25_n_489 | mul_22_25_n_355));
 assign mul_22_25_n_695 = ~((mul_22_25_n_280 | mul_22_25_n_245) & (mul_22_25_n_485 | mul_22_25_n_221));
 assign mul_22_25_n_694 = ~((mul_22_25_n_283 | mul_22_25_n_201) & (mul_22_25_n_487 | mul_22_25_n_411));
 assign mul_22_25_n_693 = ~((mul_22_25_n_287 | mul_22_25_n_224) & (mul_22_25_n_479 | mul_22_25_n_362));
 assign mul_22_25_n_692 = ~((mul_22_25_n_286 | mul_22_25_n_197) & (mul_22_25_n_483 | mul_22_25_n_290));
 assign mul_22_25_n_691 = ~((mul_22_25_n_280 | mul_22_25_n_263) & (mul_22_25_n_485 | mul_22_25_n_217));
 assign mul_22_25_n_690 = ~((mul_22_25_n_286 | mul_22_25_n_150) & (mul_22_25_n_483 | mul_22_25_n_312));
 assign mul_22_25_n_689 = ~((mul_22_25_n_284 | mul_22_25_n_107) & (mul_22_25_n_491 | mul_22_25_n_173));
 assign mul_22_25_n_688 = ~((mul_22_25_n_281 | mul_22_25_n_237) & (mul_22_25_n_493 | mul_22_25_n_264));
 assign mul_22_25_n_687 = ~((mul_22_25_n_281 | mul_22_25_n_443) & (mul_22_25_n_493 | mul_22_25_n_214));
 assign mul_22_25_n_686 = ~((mul_22_25_n_283 | mul_22_25_n_349) & (mul_22_25_n_487 | mul_22_25_n_351));
 assign mul_22_25_n_685 = ~(mul_22_25_n_505 & (mul_22_25_n_491 | mul_22_25_n_236));
 assign mul_22_25_n_684 = ~((mul_22_25_n_284 | mul_22_25_n_374) & (mul_22_25_n_491 | mul_22_25_n_291));
 assign mul_22_25_n_683 = ~((mul_22_25_n_288 | mul_22_25_n_369) & (mul_22_25_n_494 | mul_22_25_n_203));
 assign mul_22_25_n_682 = ~((mul_22_25_n_284 | mul_22_25_n_182) & (mul_22_25_n_491 | mul_22_25_n_405));
 assign mul_22_25_n_681 = ~((mul_22_25_n_280 | mul_22_25_n_393) & (mul_22_25_n_485 | mul_22_25_n_245));
 assign mul_22_25_n_680 = ~((mul_22_25_n_282 | mul_22_25_n_115) & (mul_22_25_n_481 | mul_22_25_n_114));
 assign mul_22_25_n_679 = ~((mul_22_25_n_288 | mul_22_25_n_191) & (mul_22_25_n_494 | mul_22_25_n_326));
 assign mul_22_25_n_678 = ~((mul_22_25_n_284 | mul_22_25_n_331) & (mul_22_25_n_491 | mul_22_25_n_117));
 assign mul_22_25_n_677 = ~((mul_22_25_n_287 | mul_22_25_n_110) & (mul_22_25_n_479 | mul_22_25_n_235));
 assign mul_22_25_n_676 = ~((mul_22_25_n_282 | mul_22_25_n_116) & (mul_22_25_n_481 | mul_22_25_n_188));
 assign mul_22_25_n_675 = ~((mul_22_25_n_282 | mul_22_25_n_119) & (mul_22_25_n_481 | mul_22_25_n_169));
 assign mul_22_25_n_674 = ~((mul_22_25_n_286 | mul_22_25_n_312) & (mul_22_25_n_483 | mul_22_25_n_204));
 assign mul_22_25_n_673 = ~((mul_22_25_n_287 | mul_22_25_n_365) & (mul_22_25_n_479 | mul_22_25_n_142));
 assign mul_22_25_n_672 = ~((mul_22_25_n_281 | mul_22_25_n_120) & (mul_22_25_n_493 | mul_22_25_n_443));
 assign mul_22_25_n_671 = ((mul_22_25_n_457 & mul_22_25_n_356) | (mul_22_25_n_484 & mul_22_25_n_171));
 assign mul_22_25_n_670 = ~((mul_22_25_n_287 | mul_22_25_n_422) & (mul_22_25_n_479 | mul_22_25_n_365));
 assign mul_22_25_n_669 = ~((mul_22_25_n_282 | mul_22_25_n_251) & (mul_22_25_n_481 | mul_22_25_n_115));
 assign mul_22_25_n_668 = ~((mul_22_25_n_283 | mul_22_25_n_350) & (mul_22_25_n_487 | mul_22_25_n_441));
 assign mul_22_25_n_667 = ~((mul_22_25_n_288 | mul_22_25_n_195) & (mul_22_25_n_494 | mul_22_25_n_166));
 assign mul_22_25_n_666 = ~((mul_22_25_n_282 | mul_22_25_n_169) & (mul_22_25_n_481 | mul_22_25_n_168));
 assign mul_22_25_n_665 = ~((mul_22_25_n_282 | mul_22_25_n_304) & (mul_22_25_n_481 | mul_22_25_n_156));
 assign mul_22_25_n_664 = ~((mul_22_25_n_280 | mul_22_25_n_262) & (mul_22_25_n_485 | mul_22_25_n_393));
 assign mul_22_25_n_663 = ~((mul_22_25_n_286 | mul_22_25_n_112) & (mul_22_25_n_483 | mul_22_25_n_197));
 assign mul_22_25_n_662 = ~((mul_22_25_n_284 | mul_22_25_n_405) & (mul_22_25_n_491 | mul_22_25_n_333));
 assign mul_22_25_n_661 = ~((mul_22_25_n_285 | mul_22_25_n_145) & (mul_22_25_n_489 | mul_22_25_n_364));
 assign mul_22_25_n_660 = ~((mul_22_25_n_280 | mul_22_25_n_294) & (mul_22_25_n_485 | mul_22_25_n_262));
 assign mul_22_25_n_659 = ~((mul_22_25_n_282 | mul_22_25_n_200) & (mul_22_25_n_481 | mul_22_25_n_251));
 assign mul_22_25_n_658 = ~((mul_22_25_n_285 | mul_22_25_n_109) & (mul_22_25_n_489 | mul_22_25_n_397));
 assign mul_22_25_n_657 = ~((mul_22_25_n_280 | mul_22_25_n_170) & (mul_22_25_n_485 | mul_22_25_n_294));
 assign mul_22_25_n_656 = ~((mul_22_25_n_284 | mul_22_25_n_179) & (mul_22_25_n_491 | mul_22_25_n_209));
 assign mul_22_25_n_655 = ~((mul_22_25_n_285 | mul_22_25_n_328) & (mul_22_25_n_489 | mul_22_25_n_419));
 assign mul_22_25_n_654 = ~((mul_22_25_n_284 | mul_22_25_n_415) & (mul_22_25_n_491 | mul_22_25_n_361));
 assign mul_22_25_n_653 = ~((mul_22_25_n_282 | mul_22_25_n_377) & (mul_22_25_n_481 | mul_22_25_n_119));
 assign mul_22_25_n_652 = ~((mul_22_25_n_287 | mul_22_25_n_142) & (mul_22_25_n_479 | mul_22_25_n_224));
 assign mul_22_25_n_651 = ~((mul_22_25_n_288 | mul_22_25_n_151) & (mul_22_25_n_494 | mul_22_25_n_163));
 assign mul_22_25_n_650 = ~((mul_22_25_n_282 | mul_22_25_n_188) & (mul_22_25_n_481 | mul_22_25_n_444));
 assign mul_22_25_n_649 = ~((mul_22_25_n_285 | mul_22_25_n_397) & (mul_22_25_n_489 | mul_22_25_n_292));
 assign mul_22_25_n_648 = ~((mul_22_25_n_286 | mul_22_25_n_412) & (mul_22_25_n_483 | mul_22_25_n_258));
 assign mul_22_25_n_647 = ~((mul_22_25_n_280 | mul_22_25_n_220) & (mul_22_25_n_485 | mul_22_25_n_407));
 assign mul_22_25_n_646 = ~((mul_22_25_n_287 | mul_22_25_n_389) & (mul_22_25_n_479 | mul_22_25_n_383));
 assign mul_22_25_n_645 = ~((mul_22_25_n_288 | mul_22_25_n_363) & (mul_22_25_n_494 | mul_22_25_n_386));
 assign mul_22_25_n_644 = ~((mul_22_25_n_285 | mul_22_25_n_127) & (mul_22_25_n_489 | mul_22_25_n_310));
 assign mul_22_25_n_643 = ~((mul_22_25_n_286 | mul_22_25_n_196) & (mul_22_25_n_483 | mul_22_25_n_329));
 assign mul_22_25_n_642 = ~((mul_22_25_n_287 | mul_22_25_n_244) & (mul_22_25_n_479 | mul_22_25_n_359));
 assign mul_22_25_n_641 = ~((mul_22_25_n_283 | mul_22_25_n_222) & (mul_22_25_n_487 | mul_22_25_n_350));
 assign mul_22_25_n_640 = ~((mul_22_25_n_282 | mul_22_25_n_138) & (mul_22_25_n_481 | mul_22_25_n_321));
 assign mul_22_25_n_639 = ~((mul_22_25_n_283 | mul_22_25_n_218) & (mul_22_25_n_487 | mul_22_25_n_360));
 assign mul_22_25_n_638 = ~((mul_22_25_n_282 | mul_22_25_n_325) & (mul_22_25_n_481 | mul_22_25_n_111));
 assign mul_22_25_n_637 = ~((mul_22_25_n_283 | mul_22_25_n_202) & (mul_22_25_n_487 | mul_22_25_n_222));
 assign mul_22_25_n_636 = ~((mul_22_25_n_286 | mul_22_25_n_268) & (mul_22_25_n_483 | mul_22_25_n_206));
 assign mul_22_25_n_635 = ~((mul_22_25_n_284 | mul_22_25_n_236) & (mul_22_25_n_491 | mul_22_25_n_403));
 assign mul_22_25_n_634 = ~((mul_22_25_n_282 | mul_22_25_n_212) & (mul_22_25_n_481 | mul_22_25_n_200));
 assign mul_22_25_n_633 = ~((mul_22_25_n_283 | mul_22_25_n_159) & (mul_22_25_n_487 | mul_22_25_n_201));
 assign mul_22_25_n_632 = ~((mul_22_25_n_288 | mul_22_25_n_162) & (mul_22_25_n_494 | mul_22_25_n_187));
 assign mul_22_25_n_631 = ~((mul_22_25_n_288 | mul_22_25_n_113) & (mul_22_25_n_494 | mul_22_25_n_363));
 assign mul_22_25_n_630 = ~((mul_22_25_n_287 | mul_22_25_n_184) & (mul_22_25_n_479 | mul_22_25_n_343));
 assign mul_22_25_n_629 = ~((mul_22_25_n_286 | mul_22_25_n_206) & (mul_22_25_n_483 | mul_22_25_n_136));
 assign mul_22_25_n_628 = ~((mul_22_25_n_286 | mul_22_25_n_157) & (mul_22_25_n_483 | mul_22_25_n_150));
 assign mul_22_25_n_627 = ~((mul_22_25_n_280 | mul_22_25_n_408) & (mul_22_25_n_485 | mul_22_25_n_220));
 assign mul_22_25_n_626 = ~((mul_22_25_n_285 | mul_22_25_n_160) & (mul_22_25_n_489 | mul_22_25_n_225));
 assign mul_22_25_n_625 = ~((mul_22_25_n_288 | mul_22_25_n_185) & (mul_22_25_n_494 | mul_22_25_n_398));
 assign mul_22_25_n_624 = ~((mul_22_25_n_288 | mul_22_25_n_187) & (mul_22_25_n_494 | mul_22_25_n_113));
 assign mul_22_25_n_623 = ((mul_22_25_n_454 & mul_22_25_n_427) | (mul_22_25_n_480 & mul_22_25_n_289));
 assign mul_22_25_n_622 = ~((mul_22_25_n_281 | mul_22_25_n_192) & (mul_22_25_n_493 | mul_22_25_n_165));
 assign mul_22_25_n_621 = ~((mul_22_25_n_285 | mul_22_25_n_355) & (mul_22_25_n_489 | mul_22_25_n_328));
 assign mul_22_25_n_620 = ~((mul_22_25_n_280 | mul_22_25_n_183) & (mul_22_25_n_485 | mul_22_25_n_141));
 assign mul_22_25_n_619 = ~((mul_22_25_n_286 | mul_22_25_n_372) & (mul_22_25_n_483 | mul_22_25_n_268));
 assign mul_22_25_n_618 = ~((mul_22_25_n_288 | mul_22_25_n_199) & (mul_22_25_n_494 | mul_22_25_n_158));
 assign mul_22_25_n_617 = ~((mul_22_25_n_283 | mul_22_25_n_357) & (mul_22_25_n_487 | mul_22_25_n_367));
 assign mul_22_25_n_616 = ~((mul_22_25_n_284 | mul_22_25_n_186) & (mul_22_25_n_491 | mul_22_25_n_395));
 assign mul_22_25_n_615 = ~((mul_22_25_n_284 | mul_22_25_n_442) & (mul_22_25_n_491 | mul_22_25_n_353));
 assign mul_22_25_n_614 = ~((mul_22_25_n_283 | mul_22_25_n_190) & (mul_22_25_n_487 | mul_22_25_n_381));
 assign mul_22_25_n_613 = ~((mul_22_25_n_287 | mul_22_25_n_416) & (mul_22_25_n_479 | mul_22_25_n_309));
 assign mul_22_25_n_612 = ~((mul_22_25_n_287 | mul_22_25_n_383) & (mul_22_25_n_479 | mul_22_25_n_347));
 assign mul_22_25_n_611 = ~((mul_22_25_n_284 | mul_22_25_n_209) & (mul_22_25_n_491 | mul_22_25_n_240));
 assign mul_22_25_n_610 = ~((mul_22_25_n_282 | mul_22_25_n_180) & (mul_22_25_n_481 | mul_22_25_n_448));
 assign mul_22_25_n_609 = ~((mul_22_25_n_286 | mul_22_25_n_358) & (mul_22_25_n_483 | mul_22_25_n_157));
 assign mul_22_25_n_608 = ~((mul_22_25_n_287 | mul_22_25_n_176) & (mul_22_25_n_479 | mul_22_25_n_389));
 assign mul_22_25_n_607 = ~((mul_22_25_n_288 | mul_22_25_n_388) & (mul_22_25_n_494 | mul_22_25_n_185));
 assign mul_22_25_n_606 = ~((mul_22_25_n_285 | mul_22_25_n_336) & (mul_22_25_n_489 | mul_22_25_n_160));
 assign mul_22_25_n_605 = ~((mul_22_25_n_283 | mul_22_25_n_351) & (mul_22_25_n_487 | mul_22_25_n_293));
 assign mul_22_25_n_604 = ~((mul_22_25_n_282 | mul_22_25_n_321) & (mul_22_25_n_481 | mul_22_25_n_212));
 assign mul_22_25_n_603 = ~((mul_22_25_n_280 | mul_22_25_n_228) & (mul_22_25_n_485 | mul_22_25_n_183));
 assign mul_22_25_n_602 = ~((mul_22_25_n_284 | mul_22_25_n_240) & (mul_22_25_n_491 | mul_22_25_n_311));
 assign mul_22_25_n_601 = ~((mul_22_25_n_281 | mul_22_25_n_243) & (mul_22_25_n_493 | mul_22_25_n_253));
 assign mul_22_25_n_600 = ~((mul_22_25_n_288 | mul_22_25_n_398) & (mul_22_25_n_494 | mul_22_25_n_195));
 assign mul_22_25_n_599 = ~((mul_22_25_n_288 | mul_22_25_n_386) & (mul_22_25_n_494 | mul_22_25_n_191));
 assign mul_22_25_n_598 = ~((mul_22_25_n_282 | mul_22_25_n_123) & (mul_22_25_n_481 | mul_22_25_n_198));
 assign mul_22_25_n_597 = ~((mul_22_25_n_287 | mul_22_25_n_343) & (mul_22_25_n_479 | mul_22_25_n_303));
 assign mul_22_25_n_596 = ~((mul_22_25_n_284 | mul_22_25_n_117) & (mul_22_25_n_491 | mul_22_25_n_147));
 assign mul_22_25_n_595 = ~((mul_22_25_n_283 | mul_22_25_n_367) & (mul_22_25_n_487 | mul_22_25_n_233));
 assign mul_22_25_n_594 = ~((mul_22_25_n_281 | mul_22_25_n_210) & (mul_22_25_n_493 | mul_22_25_n_192));
 assign mul_22_25_n_593 = ~((mul_22_25_n_285 | mul_22_25_n_310) & (mul_22_25_n_489 | mul_22_25_n_178));
 assign mul_22_25_n_592 = ~((mul_22_25_n_286 | mul_22_25_n_322) & (mul_22_25_n_483 | mul_22_25_n_358));
 assign mul_22_25_n_591 = ~((mul_22_25_n_285 | mul_22_25_n_152) & (mul_22_25_n_489 | mul_22_25_n_109));
 assign mul_22_25_n_590 = ~((mul_22_25_n_287 | mul_22_25_n_400) & (mul_22_25_n_479 | mul_22_25_n_176));
 assign mul_22_25_n_589 = ~((mul_22_25_n_280 | mul_22_25_n_146) & (mul_22_25_n_485 | mul_22_25_n_408));
 assign mul_22_25_n_588 = ~((mul_22_25_n_288 | mul_22_25_n_327) & (mul_22_25_n_494 | mul_22_25_n_388));
 assign mul_22_25_n_587 = ~((mul_22_25_n_280 | mul_22_25_n_149) & (mul_22_25_n_485 | mul_22_25_n_228));
 assign mul_22_25_n_586 = ~((mul_22_25_n_288 | mul_22_25_n_436) & (mul_22_25_n_494 | mul_22_25_n_121));
 assign mul_22_25_n_585 = ~((mul_22_25_n_288 | mul_22_25_n_166) & (mul_22_25_n_494 | mul_22_25_n_404));
 assign mul_22_25_n_584 = ~((mul_22_25_n_283 | mul_22_25_n_293) & (mul_22_25_n_487 | mul_22_25_n_193));
 assign mul_22_25_n_583 = ~((mul_22_25_n_280 | mul_22_25_n_227) & (mul_22_25_n_485 | mul_22_25_n_133));
 assign mul_22_25_n_582 = ~((mul_22_25_n_285 | mul_22_25_n_230) & (mul_22_25_n_489 | mul_22_25_n_302));
 assign mul_22_25_n_581 = ~((mul_22_25_n_288 | mul_22_25_n_177) & (mul_22_25_n_494 | mul_22_25_n_162));
 assign mul_22_25_n_580 = ~((mul_22_25_n_283 | mul_22_25_n_434) & (mul_22_25_n_487 | mul_22_25_n_202));
 assign mul_22_25_n_579 = ~((mul_22_25_n_285 | mul_22_25_n_178) & (mul_22_25_n_489 | mul_22_25_n_332));
 assign mul_22_25_n_578 = ~((mul_22_25_n_284 | mul_22_25_n_391) & (mul_22_25_n_491 | mul_22_25_n_374));
 assign mul_22_25_n_577 = ~((mul_22_25_n_280 | mul_22_25_n_298) & (mul_22_25_n_485 | mul_22_25_n_146));
 assign mul_22_25_n_576 = ~((mul_22_25_n_284 | mul_22_25_n_147) & (mul_22_25_n_491 | mul_22_25_n_107));
 assign mul_22_25_n_575 = ~((mul_22_25_n_284 | mul_22_25_n_361) & (mul_22_25_n_491 | mul_22_25_n_179));
 assign mul_22_25_n_574 = ~((mul_22_25_n_282 | mul_22_25_n_216) & (mul_22_25_n_481 | mul_22_25_n_123));
 assign mul_22_25_n_573 = ~((mul_22_25_n_282 | mul_22_25_n_409) & (mul_22_25_n_481 | mul_22_25_n_330));
 assign mul_22_25_n_572 = ~((mul_22_25_n_286 | mul_22_25_n_384) & (mul_22_25_n_483 | mul_22_25_n_322));
 assign mul_22_25_n_571 = ~((mul_22_25_n_287 | mul_22_25_n_122) & (mul_22_25_n_479 | mul_22_25_n_400));
 assign mul_22_25_n_570 = ~((mul_22_25_n_288 | mul_22_25_n_131) & (mul_22_25_n_494 | mul_22_25_n_327));
 assign mul_22_25_n_569 = ((mul_22_25_n_454 & mul_22_25_n_229) | (mul_22_25_n_480 & mul_22_25_n_137));
 assign mul_22_25_n_568 = ~((mul_22_25_n_281 | mul_22_25_n_256) & (mul_22_25_n_493 | mul_22_25_n_243));
 assign mul_22_25_n_567 = ~((mul_22_25_n_283 | mul_22_25_n_378) & (mul_22_25_n_487 | mul_22_25_n_349));
 assign mul_22_25_n_566 = ~((mul_22_25_n_280 | mul_22_25_n_249) & (mul_22_25_n_485 | mul_22_25_n_149));
 assign mul_22_25_n_565 = ~((mul_22_25_n_283 | mul_22_25_n_125) & (mul_22_25_n_487 | mul_22_25_n_357));
 assign mul_22_25_n_564 = ~((mul_22_25_n_283 | mul_22_25_n_181) & (mul_22_25_n_487 | mul_22_25_n_125));
 assign mul_22_25_n_563 = ~((mul_22_25_n_286 | mul_22_25_n_375) & (mul_22_25_n_483 | mul_22_25_n_412));
 assign mul_22_25_n_562 = ~((mul_22_25_n_285 | mul_22_25_n_219) & (mul_22_25_n_489 | mul_22_25_n_152));
 assign mul_22_25_n_711 = ((mul_22_25_n_284 | mul_22_25_n_353) & (mul_22_25_n_491 | mul_22_25_n_259));
 assign mul_22_25_n_710 = ~((mul_22_25_n_455 & mul_22_25_n_260) | (mul_22_25_n_492 & mul_22_25_n_205));
 assign mul_22_25_n_709 = ((mul_22_25_n_281 | mul_22_25_n_406) & (mul_22_25_n_493 | mul_22_25_n_210));
 assign mul_22_25_n_708 = ~((mul_22_25_n_455 & mul_22_25_n_205) | (mul_22_25_n_492 & mul_22_25_n_161));
 assign mul_22_25_n_707 = ((mul_22_25_n_455 & mul_22_25_n_261) | (mul_22_25_n_492 & mul_22_25_n_305));
 assign mul_22_25_n_706 = ((mul_22_25_n_455 & mul_22_25_n_154) | (mul_22_25_n_492 & mul_22_25_n_260));
 assign mul_22_25_n_705 = ~((mul_22_25_n_455 & mul_22_25_n_385) | (mul_22_25_n_492 & mul_22_25_n_261));
 assign mul_22_25_n_554 = ~((mul_22_25_n_380 | mul_22_25_n_52) & (mul_22_25_n_450 | mul_22_25_n_401));
 assign mul_22_25_n_553 = ~(({in1[18]} & {in2[0]}) | ({in1[17]} & ({in1[18]} ^ {in2[0]})));
 assign mul_22_25_n_552 = ~(({in1[2]} & {in2[0]}) | ({in1[1]} & ({in1[2]} ^ {in2[0]})));
 assign mul_22_25_n_551 = ~(({in1[8]} & {in2[0]}) | ({in1[7]} & ({in1[8]} ^ {in2[0]})));
 assign mul_22_25_n_550 = ~(({in1[10]} & {in2[0]}) | ({in1[9]} & ({in1[10]} ^ {in2[0]})));
 assign mul_22_25_n_549 = ~(({in1[6]} & {in2[0]}) | ({in1[5]} & ({in1[6]} ^ {in2[0]})));
 assign mul_22_25_n_548 = ~(({in1[14]} & {in2[0]}) | ({in1[13]} & ({in1[14]} ^ {in2[0]})));
 assign mul_22_25_n_547 = ~(({in1[12]} & {in2[0]}) | ({in1[11]} & ({in1[12]} ^ {in2[0]})));
 assign mul_22_25_n_546 = ~(({in1[16]} & {in2[0]}) | ({in1[15]} & ({in1[16]} ^ {in2[0]})));
 assign mul_22_25_n_545 = ~(({in1[4]} & {in2[0]}) | ({in1[3]} & ({in1[4]} ^ {in2[0]})));
 assign mul_22_25_n_544 = ~((mul_22_25_n_396 | mul_22_25_n_52) & (mul_22_25_n_450 | mul_22_25_n_339));
 assign mul_22_25_n_543 = ~((mul_22_25_n_306 | mul_22_25_n_52) & (mul_22_25_n_450 | mul_22_25_n_334));
 assign mul_22_25_n_561 = ~((mul_22_25_n_118 & {in1[0]}) | (mul_22_25_n_451 & mul_22_25_n_94));
 assign mul_22_25_n_560 = ~((mul_22_25_n_108 & {in1[0]}) | (mul_22_25_n_451 & mul_22_25_n_213));
 assign mul_22_25_n_559 = ~(mul_22_25_n_452 & (mul_22_25_n_450 | mul_22_25_n_421));
 assign mul_22_25_n_558 = ~((mul_22_25_n_269 & {in1[0]}) | (mul_22_25_n_451 & mul_22_25_n_108));
 assign mul_22_25_n_557 = ~((mul_22_25_n_340 & {in1[0]}) | (mul_22_25_n_451 & mul_22_25_n_307));
 assign mul_22_25_n_556 = ~((mul_22_25_n_194 & {in1[0]}) | (mul_22_25_n_451 & mul_22_25_n_269));
 assign mul_22_25_n_555 = ~((mul_22_25_n_342 & {in1[0]}) | (mul_22_25_n_451 & mul_22_25_n_172));
 assign mul_22_25_n_530 = ((mul_22_25_n_172 & {in1[0]}) | (mul_22_25_n_451 & mul_22_25_n_323));
 assign mul_22_25_n_529 = ~((mul_22_25_n_320 | mul_22_25_n_52) & (mul_22_25_n_450 | mul_22_25_n_440));
 assign mul_22_25_n_528 = ~((mul_22_25_n_167 | mul_22_25_n_52) & (mul_22_25_n_450 | mul_22_25_n_380));
 assign mul_22_25_n_527 = ~((mul_22_25_n_401 | mul_22_25_n_52) & (mul_22_25_n_450 | mul_22_25_n_132));
 assign mul_22_25_n_526 = ~((mul_22_25_n_300 | mul_22_25_n_52) & (mul_22_25_n_450 | mul_22_25_n_315));
 assign mul_22_25_n_525 = ~((mul_22_25_n_132 | mul_22_25_n_52) & (mul_22_25_n_450 | mul_22_25_n_345));
 assign mul_22_25_n_524 = ((mul_22_25_n_153 & {in1[0]}) | (mul_22_25_n_451 & mul_22_25_n_342));
 assign mul_22_25_n_523 = ~(mul_22_25_n_449 & (mul_22_25_n_450 | mul_22_25_n_396));
 assign mul_22_25_n_522 = ~((mul_22_25_n_128 | mul_22_25_n_52) & (mul_22_25_n_450 | mul_22_25_n_167));
 assign mul_22_25_n_542 = ~((mul_22_25_n_297 & {in1[0]}) | (mul_22_25_n_451 & mul_22_25_n_118));
 assign mul_22_25_n_541 = ~((mul_22_25_n_346 & {in1[0]}) | (mul_22_25_n_451 & mul_22_25_n_301));
 assign mul_22_25_n_540 = ~((~mul_22_25_n_334 & ~mul_22_25_n_52) | (mul_22_25_n_451 & mul_22_25_n_153));
 assign mul_22_25_n_539 = ~((mul_22_25_n_134 & {in1[0]}) | (mul_22_25_n_451 & mul_22_25_n_194));
 assign mul_22_25_n_538 = ~((~mul_22_25_n_421 & ~mul_22_25_n_52) | (mul_22_25_n_451 & mul_22_25_n_140));
 assign mul_22_25_n_537 = ~((mul_22_25_n_439 & {in1[0]}) | (mul_22_25_n_451 & mul_22_25_n_297));
 assign mul_22_25_n_536 = ~((mul_22_25_n_234 & {in1[0]}) | (mul_22_25_n_451 & mul_22_25_n_134));
 assign mul_22_25_n_535 = ~((mul_22_25_n_208 & {in1[0]}) | (mul_22_25_n_451 & mul_22_25_n_239));
 assign mul_22_25_n_534 = ~((mul_22_25_n_239 & {in1[0]}) | (mul_22_25_n_451 & mul_22_25_n_234));
 assign mul_22_25_n_533 = ~((mul_22_25_n_140 & {in1[0]}) | (mul_22_25_n_451 & mul_22_25_n_208));
 assign mul_22_25_n_532 = ~((mul_22_25_n_316 & {in1[0]}) | (mul_22_25_n_451 & mul_22_25_n_319));
 assign mul_22_25_n_531 = ~((mul_22_25_n_323 & {in1[0]}) | (mul_22_25_n_451 & mul_22_25_n_129));
 assign mul_22_25_n_519 = ~mul_22_25_n_2;
 assign mul_22_25_n_518 = ~mul_22_25_n_4;
 assign mul_22_25_n_514 = ~(mul_22_25_n_105 | mul_22_25_n_23);
 assign mul_22_25_n_513 = ~(mul_22_25_n_285 | mul_22_25_n_23);
 assign mul_22_25_n_512 = ~(mul_22_25_n_288 | mul_22_25_n_23);
 assign mul_22_25_n_511 = ~(mul_22_25_n_283 | mul_22_25_n_23);
 assign mul_22_25_n_510 = ~(mul_22_25_n_284 | mul_22_25_n_23);
 assign mul_22_25_n_509 = ~(mul_22_25_n_280 | mul_22_25_n_23);
 assign mul_22_25_n_508 = ~(mul_22_25_n_287 | mul_22_25_n_23);
 assign mul_22_25_n_507 = ~(mul_22_25_n_286 | mul_22_25_n_23);
 assign mul_22_25_n_506 = ~(mul_22_25_n_282 | mul_22_25_n_23);
 assign mul_22_25_n_505 = ~(mul_22_25_n_456 & mul_22_25_n_428);
 assign mul_22_25_n_504 = ~(mul_22_25_n_105 | (mul_22_25_n_70 & ({in2[6]} | mul_22_25_n_51)));
 assign mul_22_25_n_503 = ~(mul_22_25_n_105 | (mul_22_25_n_71 & ({in2[9]} | mul_22_25_n_51)));
 assign mul_22_25_n_502 = ~(mul_22_25_n_105 | (mul_22_25_n_76 & ({in2[10]} | mul_22_25_n_51)));
 assign mul_22_25_n_501 = ~(mul_22_25_n_105 | (mul_22_25_n_68 & ({in2[4]} | mul_22_25_n_51)));
 assign mul_22_25_n_500 = ~(mul_22_25_n_105 | (mul_22_25_n_67 & ({in2[21]} | mul_22_25_n_51)));
 assign mul_22_25_n_499 = ~(mul_22_25_n_105 | (mul_22_25_n_88 & ({in2[28]} | mul_22_25_n_51)));
 assign mul_22_25_n_498 = ~(mul_22_25_n_105 | (mul_22_25_n_85 & ({in2[11]} | mul_22_25_n_51)));
 assign mul_22_25_n_497 = ~(mul_22_25_n_105 | (mul_22_25_n_65 & ({in2[13]} | mul_22_25_n_51)));
 assign mul_22_25_n_496 = ~(mul_22_25_n_105 | (mul_22_25_n_91 & ({in2[12]} | mul_22_25_n_51)));
 assign mul_22_25_n_495 = ~(mul_22_25_n_105 | (mul_22_25_n_77 & ({in2[3]} | mul_22_25_n_51)));
 assign mul_22_25_n_521 = ~(mul_22_25_n_457 & mul_22_25_n_435);
 assign mul_22_25_n_520 = (mul_22_25_n_456 & mul_22_25_n_438);
 assign mul_22_25_n_517 = ~(mul_22_25_n_455 & mul_22_25_n_424);
 assign mul_22_25_n_516 = ~(mul_22_25_n_455 & {in2[0]});
 assign mul_22_25_n_515 = (mul_22_25_n_454 & mul_22_25_n_420);
 assign mul_22_25_n_492 = ~mul_22_25_n_493;
 assign mul_22_25_n_490 = ~mul_22_25_n_491;
 assign mul_22_25_n_488 = ~mul_22_25_n_489;
 assign mul_22_25_n_486 = ~mul_22_25_n_487;
 assign mul_22_25_n_484 = ~mul_22_25_n_485;
 assign mul_22_25_n_482 = ~mul_22_25_n_483;
 assign mul_22_25_n_480 = ~mul_22_25_n_481;
 assign mul_22_25_n_478 = ~mul_22_25_n_479;
 assign mul_22_25_n_477 = ~(mul_22_25_n_105 | (mul_22_25_n_81 & ({in2[5]} | mul_22_25_n_51)));
 assign mul_22_25_n_476 = ~(mul_22_25_n_105 | (mul_22_25_n_83 & ({in2[8]} | mul_22_25_n_51)));
 assign mul_22_25_n_475 = ~(mul_22_25_n_105 | (mul_22_25_n_73 & ({in2[16]} | mul_22_25_n_51)));
 assign mul_22_25_n_474 = ~(mul_22_25_n_105 | (mul_22_25_n_66 & ({in2[24]} | mul_22_25_n_51)));
 assign mul_22_25_n_473 = ~(mul_22_25_n_105 | (mul_22_25_n_80 & ({in2[2]} | mul_22_25_n_51)));
 assign mul_22_25_n_472 = ~(mul_22_25_n_105 | (mul_22_25_n_86 & ({in2[27]} | mul_22_25_n_51)));
 assign mul_22_25_n_471 = ~(mul_22_25_n_105 | (mul_22_25_n_69 & ({in2[18]} | mul_22_25_n_51)));
 assign mul_22_25_n_470 = ~(mul_22_25_n_105 | (mul_22_25_n_75 & ({in2[17]} | mul_22_25_n_51)));
 assign mul_22_25_n_469 = ~(mul_22_25_n_453 & (mul_22_25_n_74 | (mul_22_25_n_51 & {in2[29]})));
 assign mul_22_25_n_468 = ~(mul_22_25_n_105 | (mul_22_25_n_64 & ({in2[25]} | mul_22_25_n_51)));
 assign mul_22_25_n_467 = ~(mul_22_25_n_105 | (mul_22_25_n_82 & ({in2[15]} | mul_22_25_n_51)));
 assign mul_22_25_n_466 = ~(mul_22_25_n_105 | (mul_22_25_n_90 & ({in2[26]} | mul_22_25_n_51)));
 assign mul_22_25_n_465 = ~(mul_22_25_n_105 | (mul_22_25_n_92 & ({in2[19]} | mul_22_25_n_51)));
 assign mul_22_25_n_464 = ~(mul_22_25_n_105 | (mul_22_25_n_78 & ({in2[22]} | mul_22_25_n_51)));
 assign mul_22_25_n_463 = ~(mul_22_25_n_105 | (mul_22_25_n_87 & ({in2[14]} | mul_22_25_n_51)));
 assign mul_22_25_n_462 = ~(mul_22_25_n_105 | (mul_22_25_n_79 & ({in2[23]} | mul_22_25_n_51)));
 assign mul_22_25_n_461 = ~(mul_22_25_n_105 | (mul_22_25_n_72 & ({in2[1]} | mul_22_25_n_51)));
 assign mul_22_25_n_460 = ~(mul_22_25_n_105 | (mul_22_25_n_84 & ({in2[7]} | mul_22_25_n_51)));
 assign mul_22_25_n_459 = ~(mul_22_25_n_105 | (mul_22_25_n_89 & ({in2[20]} | mul_22_25_n_51)));
 assign mul_22_25_n_494 = ~(mul_22_25_n_288 & mul_22_25_n_278);
 assign mul_22_25_n_493 = ~(mul_22_25_n_281 & mul_22_25_n_272);
 assign mul_22_25_n_491 = ~(mul_22_25_n_284 & mul_22_25_n_276);
 assign mul_22_25_n_489 = ~(mul_22_25_n_285 & mul_22_25_n_275);
 assign mul_22_25_n_487 = ~(mul_22_25_n_283 & mul_22_25_n_279);
 assign mul_22_25_n_485 = ~(mul_22_25_n_280 & mul_22_25_n_277);
 assign mul_22_25_n_483 = ~(mul_22_25_n_286 & mul_22_25_n_274);
 assign mul_22_25_n_481 = ~(mul_22_25_n_282 & mul_22_25_n_273);
 assign mul_22_25_n_479 = ~(mul_22_25_n_287 & mul_22_25_n_271);
 assign mul_22_25_n_457 = ~mul_22_25_n_280;
 assign mul_22_25_n_456 = ~mul_22_25_n_284;
 assign mul_22_25_n_455 = ~mul_22_25_n_281;
 assign mul_22_25_n_454 = ~mul_22_25_n_282;
 assign mul_22_25_n_453 = ~mul_22_25_n_105;
 assign mul_22_25_n_452 = ~(mul_22_25_n_430 & {in1[0]});
 assign mul_22_25_n_450 = ~mul_22_25_n_451;
 assign mul_22_25_n_449 = ~(mul_22_25_n_213 & {in1[0]});
 assign mul_22_25_n_451 = ~(mul_22_25_n_44 | {in1[0]});
 assign mul_22_25_n_440 = ~mul_22_25_n_439;
 assign mul_22_25_n_433 = ~mul_22_25_n_432;
 assign mul_22_25_n_426 = ~mul_22_25_n_425;
 assign mul_22_25_n_346 = ~mul_22_25_n_345;
 assign mul_22_25_n_340 = ~mul_22_25_n_339;
 assign mul_22_25_n_320 = ~mul_22_25_n_319;
 assign mul_22_25_n_316 = ~mul_22_25_n_315;
 assign mul_22_25_n_307 = ~mul_22_25_n_306;
 assign mul_22_25_n_301 = ~mul_22_25_n_300;
 assign mul_22_25_n_279 = ~((mul_22_25_n_49 & ~{in1[10]}) | ({in1[11]} & {in1[10]}));
 assign mul_22_25_n_278 = ~((mul_22_25_n_45 & ~{in1[18]}) | ({in1[19]} & {in1[18]}));
 assign mul_22_25_n_277 = ~((mul_22_25_n_21 & ~{in1[12]}) | ({in1[13]} & {in1[12]}));
 assign mul_22_25_n_276 = ~((mul_22_25_n_48 & ~{in1[6]}) | ({in1[7]} & {in1[6]}));
 assign mul_22_25_n_275 = ~((mul_22_25_n_20 & ~{in1[4]}) | ({in1[5]} & {in1[4]}));
 assign mul_22_25_n_274 = ~((mul_22_25_n_22 & ~{in1[16]}) | ({in1[17]} & {in1[16]}));
 assign mul_22_25_n_273 = ~((mul_22_25_n_50 & ~{in1[14]}) | ({in1[15]} & {in1[14]}));
 assign mul_22_25_n_272 = ~((mul_22_25_n_47 & ~{in1[2]}) | ({in1[3]} & {in1[2]}));
 assign mul_22_25_n_271 = ~((mul_22_25_n_46 & ~{in1[8]}) | ({in1[9]} & {in1[8]}));
 assign mul_22_25_n_270 = ~((mul_22_25_n_42 & {in1[19]}) | (mul_22_25_n_45 & {in2[31]}));
 assign mul_22_25_n_448 = ~((mul_22_25_n_37 & {in1[15]}) | (mul_22_25_n_50 & {in2[10]}));
 assign mul_22_25_n_447 = ~({in1[1]} & ~asc001_0_);
 assign mul_22_25_n_446 = ~((mul_22_25_n_41 & {in1[17]}) | (mul_22_25_n_22 & {in2[13]}));
 assign mul_22_25_n_445 = ~((mul_22_25_n_37 & {in1[3]}) | (mul_22_25_n_47 & {in2[10]}));
 assign mul_22_25_n_444 = ~((mul_22_25_n_30 & {in1[15]}) | (mul_22_25_n_50 & {in2[18]}));
 assign mul_22_25_n_443 = ~((mul_22_25_n_29 & {in1[3]}) | (mul_22_25_n_47 & {in2[2]}));
 assign mul_22_25_n_442 = ~((mul_22_25_n_57 & {in1[7]}) | (mul_22_25_n_48 & {in2[27]}));
 assign mul_22_25_n_441 = ~((mul_22_25_n_24 & {in1[11]}) | (mul_22_25_n_49 & {in2[26]}));
 assign mul_22_25_n_439 = ~(({in2[3]} | mul_22_25_n_44) & ({in1[1]} | mul_22_25_n_58));
 assign mul_22_25_n_438 = ~(({in2[31]} | mul_22_25_n_48) & ({in1[7]} | mul_22_25_n_42));
 assign mul_22_25_n_437 = ~((mul_22_25_n_43 & {in1[13]}) | (mul_22_25_n_21 & {in2[30]}));
 assign mul_22_25_n_436 = ~((mul_22_25_n_43 & {in1[19]}) | (mul_22_25_n_45 & {in2[30]}));
 assign mul_22_25_n_435 = ~(({in2[31]} | mul_22_25_n_21) & ({in1[13]} | mul_22_25_n_42));
 assign mul_22_25_n_434 = ~((mul_22_25_n_43 & {in1[11]}) | (mul_22_25_n_49 & {in2[30]}));
 assign mul_22_25_n_432 = ~(({in2[30]} | mul_22_25_n_22) & ({in1[17]} | mul_22_25_n_43));
 assign mul_22_25_n_431 = ~(({in2[31]} | mul_22_25_n_46) & ({in1[9]} | mul_22_25_n_42));
 assign mul_22_25_n_430 = ~(({in2[31]} | mul_22_25_n_44) & ({in1[1]} | mul_22_25_n_42));
 assign mul_22_25_n_429 = ~(({in2[31]} | mul_22_25_n_20) & ({in1[5]} | mul_22_25_n_42));
 assign mul_22_25_n_428 = ~(({in2[30]} | mul_22_25_n_48) & ({in1[7]} | mul_22_25_n_43));
 assign mul_22_25_n_427 = ~(({in2[30]} | mul_22_25_n_50) & ({in1[15]} | mul_22_25_n_43));
 assign mul_22_25_n_425 = ~((mul_22_25_n_43 & {in1[3]}) | (mul_22_25_n_47 & {in2[30]}));
 assign mul_22_25_n_424 = ~(({in2[31]} | mul_22_25_n_47) & ({in1[3]} | mul_22_25_n_42));
 assign mul_22_25_n_423 = ~((mul_22_25_n_43 & {in1[5]}) | (mul_22_25_n_20 & {in2[30]}));
 assign mul_22_25_n_422 = ~((mul_22_25_n_43 & {in1[9]}) | (mul_22_25_n_46 & {in2[30]}));
 assign mul_22_25_n_421 = ~((mul_22_25_n_43 & {in1[1]}) | (mul_22_25_n_44 & {in2[30]}));
 assign mul_22_25_n_420 = ~(({in2[31]} | mul_22_25_n_50) & ({in1[15]} | mul_22_25_n_42));
 assign mul_22_25_n_419 = ~((mul_22_25_n_36 & {in1[5]}) | (mul_22_25_n_20 & {in2[14]}));
 assign mul_22_25_n_418 = ~(({in2[31]} | mul_22_25_n_49) & ({in1[11]} | mul_22_25_n_42));
 assign mul_22_25_n_417 = ~(({in2[31]} | mul_22_25_n_22) & ({in1[17]} | mul_22_25_n_42));
 assign mul_22_25_n_416 = ~((mul_22_25_n_63 & {in1[9]}) | (mul_22_25_n_46 & {in2[6]}));
 assign mul_22_25_n_415 = ~((mul_22_25_n_61 & {in1[7]}) | (mul_22_25_n_48 & {in2[22]}));
 assign mul_22_25_n_414 = ~((mul_22_25_n_26 & {in1[17]}) | (mul_22_25_n_22 & {in2[12]}));
 assign mul_22_25_n_413 = ~((mul_22_25_n_37 & {in1[13]}) | (mul_22_25_n_21 & {in2[10]}));
 assign mul_22_25_n_412 = ~((mul_22_25_n_59 & {in1[17]}) | (mul_22_25_n_22 & {in2[24]}));
 assign mul_22_25_n_411 = ~((mul_22_25_n_37 & {in1[11]}) | (mul_22_25_n_49 & {in2[10]}));
 assign mul_22_25_n_410 = ~((mul_22_25_n_54 & {in1[17]}) | (mul_22_25_n_22 & {in2[21]}));
 assign mul_22_25_n_409 = ~((mul_22_25_n_41 & {in1[15]}) | (mul_22_25_n_50 & {in2[13]}));
 assign mul_22_25_n_408 = ~((mul_22_25_n_58 & {in1[13]}) | (mul_22_25_n_21 & {in2[3]}));
 assign mul_22_25_n_407 = ~((mul_22_25_n_38 & {in1[13]}) | (mul_22_25_n_21 & {in2[1]}));
 assign mul_22_25_n_406 = ~((mul_22_25_n_35 & {in1[3]}) | (mul_22_25_n_47 & {in2[7]}));
 assign mul_22_25_n_405 = ~((mul_22_25_n_35 & {in1[7]}) | (mul_22_25_n_48 & {in2[7]}));
 assign mul_22_25_n_404 = ~((mul_22_25_n_29 & {in1[19]}) | (mul_22_25_n_45 & {in2[2]}));
 assign mul_22_25_n_403 = ~((mul_22_25_n_39 & {in1[7]}) | (mul_22_25_n_48 & {in2[28]}));
 assign mul_22_25_n_402 = ~((mul_22_25_n_28 & {in1[9]}) | (mul_22_25_n_46 & {in2[25]}));
 assign mul_22_25_n_401 = ~((mul_22_25_n_31 & {in1[1]}) | (mul_22_25_n_44 & {in2[9]}));
 assign mul_22_25_n_400 = ~((mul_22_25_n_30 & {in1[9]}) | (mul_22_25_n_46 & {in2[18]}));
 assign mul_22_25_n_399 = ~((mul_22_25_n_63 & {in1[5]}) | (mul_22_25_n_20 & {in2[6]}));
 assign mul_22_25_n_398 = ~((mul_22_25_n_56 & {in1[19]}) | (mul_22_25_n_45 & {in2[5]}));
 assign mul_22_25_n_397 = ~((mul_22_25_n_29 & {in1[5]}) | (mul_22_25_n_20 & {in2[2]}));
 assign mul_22_25_n_396 = ~((mul_22_25_n_55 & {in1[1]}) | (mul_22_25_n_44 & {in2[20]}));
 assign mul_22_25_n_395 = ~((mul_22_25_n_25 & {in1[7]}) | (mul_22_25_n_48 & {in2[4]}));
 assign mul_22_25_n_394 = ~((mul_22_25_n_34 & {in1[11]}) | (mul_22_25_n_49 & {in2[19]}));
 assign mul_22_25_n_393 = ~((mul_22_25_n_59 & {in1[13]}) | (mul_22_25_n_21 & {in2[24]}));
 assign mul_22_25_n_392 = ~((mul_22_25_n_41 & {in1[19]}) | (mul_22_25_n_45 & {in2[13]}));
 assign mul_22_25_n_391 = ~((mul_22_25_n_58 & {in1[7]}) | (mul_22_25_n_48 & {in2[3]}));
 assign mul_22_25_n_390 = ~((mul_22_25_n_26 & {in1[3]}) | (mul_22_25_n_47 & {in2[12]}));
 assign mul_22_25_n_389 = ~((mul_22_25_n_27 & {in1[9]}) | (mul_22_25_n_46 & {in2[16]}));
 assign mul_22_25_n_388 = ~((mul_22_25_n_35 & {in1[19]}) | (mul_22_25_n_45 & {in2[7]}));
 assign mul_22_25_n_387 = ~((mul_22_25_n_32 & {in1[3]}) | (mul_22_25_n_47 & {in2[8]}));
 assign mul_22_25_n_386 = ~((mul_22_25_n_60 & {in1[19]}) | (mul_22_25_n_45 & {in2[23]}));
 assign mul_22_25_n_385 = ~(({in2[21]} | mul_22_25_n_47) & ({in1[3]} | mul_22_25_n_54));
 assign mul_22_25_n_384 = ~((mul_22_25_n_62 & {in1[17]}) | (mul_22_25_n_22 & {in2[11]}));
 assign mul_22_25_n_383 = ~((mul_22_25_n_40 & {in1[9]}) | (mul_22_25_n_46 & {in2[15]}));
 assign mul_22_25_n_382 = ~((mul_22_25_n_25 & {in1[17]}) | (mul_22_25_n_22 & {in2[4]}));
 assign mul_22_25_n_381 = ~((mul_22_25_n_59 & {in1[11]}) | (mul_22_25_n_49 & {in2[24]}));
 assign mul_22_25_n_380 = ~((mul_22_25_n_37 & {in1[1]}) | (mul_22_25_n_44 & {in2[10]}));
 assign mul_22_25_n_379 = ~((mul_22_25_n_27 & {in1[13]}) | (mul_22_25_n_21 & {in2[16]}));
 assign mul_22_25_n_378 = ~((mul_22_25_n_33 & {in1[11]}) | (mul_22_25_n_49 & {in2[17]}));
 assign mul_22_25_n_377 = ~((mul_22_25_n_31 & {in1[15]}) | (mul_22_25_n_50 & {in2[9]}));
 assign mul_22_25_n_376 = ~((mul_22_25_n_54 & {in1[13]}) | (mul_22_25_n_21 & {in2[21]}));
 assign mul_22_25_n_375 = ~((mul_22_25_n_28 & {in1[17]}) | (mul_22_25_n_22 & {in2[25]}));
 assign mul_22_25_n_374 = ~((mul_22_25_n_29 & {in1[7]}) | (mul_22_25_n_48 & {in2[2]}));
 assign mul_22_25_n_373 = ~((mul_22_25_n_28 & {in1[5]}) | (mul_22_25_n_20 & {in2[25]}));
 assign mul_22_25_n_372 = ~((mul_22_25_n_53 & {in1[17]}) | (mul_22_25_n_22 & {in2[29]}));
 assign mul_22_25_n_371 = ~((mul_22_25_n_61 & {in1[11]}) | (mul_22_25_n_49 & {in2[22]}));
 assign mul_22_25_n_370 = ~((mul_22_25_n_26 & {in1[19]}) | (mul_22_25_n_45 & {in2[12]}));
 assign mul_22_25_n_369 = ~((mul_22_25_n_30 & {in1[19]}) | (mul_22_25_n_45 & {in2[18]}));
 assign mul_22_25_n_368 = ~((mul_22_25_n_34 & {in1[13]}) | (mul_22_25_n_21 & {in2[19]}));
 assign mul_22_25_n_367 = ~((mul_22_25_n_25 & {in1[11]}) | (mul_22_25_n_49 & {in2[4]}));
 assign mul_22_25_n_366 = ~((mul_22_25_n_60 & {in1[11]}) | (mul_22_25_n_49 & {in2[23]}));
 assign mul_22_25_n_365 = ~((mul_22_25_n_53 & {in1[9]}) | (mul_22_25_n_46 & {in2[29]}));
 assign mul_22_25_n_364 = ~((mul_22_25_n_34 & {in1[5]}) | (mul_22_25_n_20 & {in2[19]}));
 assign mul_22_25_n_363 = ~((mul_22_25_n_59 & {in1[19]}) | (mul_22_25_n_45 & {in2[24]}));
 assign mul_22_25_n_362 = ~((mul_22_25_n_24 & {in1[9]}) | (mul_22_25_n_46 & {in2[26]}));
 assign mul_22_25_n_361 = ~((mul_22_25_n_54 & {in1[7]}) | (mul_22_25_n_48 & {in2[21]}));
 assign mul_22_25_n_360 = ~((mul_22_25_n_55 & {in1[11]}) | (mul_22_25_n_49 & {in2[20]}));
 assign mul_22_25_n_359 = ~((mul_22_25_n_29 & {in1[9]}) | (mul_22_25_n_46 & {in2[2]}));
 assign mul_22_25_n_358 = ~((mul_22_25_n_31 & {in1[17]}) | (mul_22_25_n_22 & {in2[9]}));
 assign mul_22_25_n_357 = ~((mul_22_25_n_56 & {in1[11]}) | (mul_22_25_n_49 & {in2[5]}));
 assign mul_22_25_n_356 = ~(({in2[28]} | mul_22_25_n_21) & ({in1[13]} | mul_22_25_n_39));
 assign mul_22_25_n_355 = ~((mul_22_25_n_27 & {in1[5]}) | (mul_22_25_n_20 & {in2[16]}));
 assign mul_22_25_n_354 = ~((mul_22_25_n_54 & {in1[9]}) | (mul_22_25_n_46 & {in2[21]}));
 assign mul_22_25_n_353 = ~((mul_22_25_n_24 & {in1[7]}) | (mul_22_25_n_48 & {in2[26]}));
 assign mul_22_25_n_352 = ~((mul_22_25_n_37 & {in1[9]}) | (mul_22_25_n_46 & {in2[10]}));
 assign mul_22_25_n_351 = ~((mul_22_25_n_40 & {in1[11]}) | (mul_22_25_n_49 & {in2[15]}));
 assign mul_22_25_n_350 = ~((mul_22_25_n_57 & {in1[11]}) | (mul_22_25_n_49 & {in2[27]}));
 assign mul_22_25_n_349 = ~((mul_22_25_n_27 & {in1[11]}) | (mul_22_25_n_49 & {in2[16]}));
 assign mul_22_25_n_348 = ~((mul_22_25_n_62 & {in1[19]}) | (mul_22_25_n_45 & {in2[11]}));
 assign mul_22_25_n_347 = ~((mul_22_25_n_36 & {in1[9]}) | (mul_22_25_n_46 & {in2[14]}));
 assign mul_22_25_n_345 = ~((mul_22_25_n_35 & {in1[1]}) | (mul_22_25_n_44 & {in2[7]}));
 assign mul_22_25_n_344 = ~((mul_22_25_n_31 & {in1[11]}) | (mul_22_25_n_49 & {in2[9]}));
 assign mul_22_25_n_343 = ~((mul_22_25_n_32 & {in1[9]}) | (mul_22_25_n_46 & {in2[8]}));
 assign mul_22_25_n_342 = ~(({in2[15]} | mul_22_25_n_44) & ({in1[1]} | mul_22_25_n_40));
 assign mul_22_25_n_341 = ~(({in2[29]} | mul_22_25_n_47) & ({in1[3]} | mul_22_25_n_53));
 assign mul_22_25_n_339 = ~((mul_22_25_n_34 & {in1[1]}) | (mul_22_25_n_44 & {in2[19]}));
 assign mul_22_25_n_338 = ~((mul_22_25_n_62 & {in1[9]}) | (mul_22_25_n_46 & {in2[11]}));
 assign mul_22_25_n_337 = ~((mul_22_25_n_36 & {in1[15]}) | (mul_22_25_n_50 & {in2[14]}));
 assign mul_22_25_n_336 = ~((mul_22_25_n_60 & {in1[5]}) | (mul_22_25_n_20 & {in2[23]}));
 assign mul_22_25_n_335 = ~((mul_22_25_n_59 & {in1[7]}) | (mul_22_25_n_48 & {in2[24]}));
 assign mul_22_25_n_334 = ~((mul_22_25_n_33 & {in1[1]}) | (mul_22_25_n_44 & {in2[17]}));
 assign mul_22_25_n_333 = ~((mul_22_25_n_63 & {in1[7]}) | (mul_22_25_n_48 & {in2[6]}));
 assign mul_22_25_n_332 = ~((mul_22_25_n_37 & {in1[5]}) | (mul_22_25_n_20 & {in2[10]}));
 assign mul_22_25_n_331 = ~((mul_22_25_n_27 & {in1[7]}) | (mul_22_25_n_48 & {in2[16]}));
 assign mul_22_25_n_330 = ~((mul_22_25_n_26 & {in1[15]}) | (mul_22_25_n_50 & {in2[12]}));
 assign mul_22_25_n_329 = ~((mul_22_25_n_29 & {in1[17]}) | (mul_22_25_n_22 & {in2[2]}));
 assign mul_22_25_n_328 = ~((mul_22_25_n_40 & {in1[5]}) | (mul_22_25_n_20 & {in2[15]}));
 assign mul_22_25_n_327 = ~((mul_22_25_n_32 & {in1[19]}) | (mul_22_25_n_45 & {in2[8]}));
 assign mul_22_25_n_326 = ~((mul_22_25_n_54 & {in1[19]}) | (mul_22_25_n_45 & {in2[21]}));
 assign mul_22_25_n_325 = ~((mul_22_25_n_56 & {in1[15]}) | (mul_22_25_n_50 & {in2[5]}));
 assign mul_22_25_n_324 = ~((mul_22_25_n_39 & {in1[5]}) | (mul_22_25_n_20 & {in2[28]}));
 assign mul_22_25_n_323 = ~(({in2[13]} | mul_22_25_n_44) & ({in1[1]} | mul_22_25_n_41));
 assign mul_22_25_n_322 = ~((mul_22_25_n_37 & {in1[17]}) | (mul_22_25_n_22 & {in2[10]}));
 assign mul_22_25_n_321 = ~((mul_22_25_n_24 & {in1[15]}) | (mul_22_25_n_50 & {in2[26]}));
 assign mul_22_25_n_319 = ~(({in2[4]} | mul_22_25_n_44) & ({in1[1]} | mul_22_25_n_25));
 assign mul_22_25_n_318 = ~((mul_22_25_n_60 & {in1[7]}) | (mul_22_25_n_48 & {in2[23]}));
 assign mul_22_25_n_317 = ~((mul_22_25_n_38 & {in1[17]}) | (mul_22_25_n_22 & {in2[1]}));
 assign mul_22_25_n_315 = ~((mul_22_25_n_56 & {in1[1]}) | (mul_22_25_n_44 & {in2[5]}));
 assign mul_22_25_n_314 = ~((mul_22_25_n_30 & {in1[5]}) | (mul_22_25_n_20 & {in2[18]}));
 assign mul_22_25_n_313 = ~((mul_22_25_n_40 & {in1[15]}) | (mul_22_25_n_50 & {in2[15]}));
 assign mul_22_25_n_312 = ~((mul_22_25_n_63 & {in1[17]}) | (mul_22_25_n_22 & {in2[6]}));
 assign mul_22_25_n_311 = ~((mul_22_25_n_33 & {in1[7]}) | (mul_22_25_n_48 & {in2[17]}));
 assign mul_22_25_n_310 = ~((mul_22_25_n_26 & {in1[5]}) | (mul_22_25_n_20 & {in2[12]}));
 assign mul_22_25_n_309 = ~((mul_22_25_n_56 & {in1[9]}) | (mul_22_25_n_46 & {in2[5]}));
 assign mul_22_25_n_308 = ~((mul_22_25_n_61 & {in1[17]}) | (mul_22_25_n_22 & {in2[22]}));
 assign mul_22_25_n_306 = ~((mul_22_25_n_30 & {in1[1]}) | (mul_22_25_n_44 & {in2[18]}));
 assign mul_22_25_n_305 = ~(({in2[19]} | mul_22_25_n_47) & ({in1[3]} | mul_22_25_n_34));
 assign mul_22_25_n_304 = ~((mul_22_25_n_33 & {in1[15]}) | (mul_22_25_n_50 & {in2[17]}));
 assign mul_22_25_n_303 = ~((mul_22_25_n_35 & {in1[9]}) | (mul_22_25_n_46 & {in2[7]}));
 assign mul_22_25_n_302 = ~((mul_22_25_n_32 & {in1[5]}) | (mul_22_25_n_20 & {in2[8]}));
 assign mul_22_25_n_300 = ~((mul_22_25_n_63 & {in1[1]}) | (mul_22_25_n_44 & {in2[6]}));
 assign mul_22_25_n_299 = ~((mul_22_25_n_62 & {in1[3]}) | (mul_22_25_n_47 & {in2[11]}));
 assign mul_22_25_n_298 = ~((mul_22_25_n_56 & {in1[13]}) | (mul_22_25_n_21 & {in2[5]}));
 assign mul_22_25_n_297 = ~(({in2[2]} | mul_22_25_n_44) & ({in1[1]} | mul_22_25_n_29));
 assign mul_22_25_n_296 = ~((mul_22_25_n_33 & {in1[13]}) | (mul_22_25_n_21 & {in2[17]}));
 assign mul_22_25_n_295 = ~((mul_22_25_n_36 & {in1[19]}) | (mul_22_25_n_45 & {in2[14]}));
 assign mul_22_25_n_294 = ~((mul_22_25_n_24 & {in1[13]}) | (mul_22_25_n_21 & {in2[26]}));
 assign mul_22_25_n_293 = ~((mul_22_25_n_36 & {in1[11]}) | (mul_22_25_n_49 & {in2[14]}));
 assign mul_22_25_n_292 = ~((mul_22_25_n_38 & {in1[5]}) | (mul_22_25_n_20 & {in2[1]}));
 assign mul_22_25_n_291 = ~((mul_22_25_n_38 & {in1[7]}) | (mul_22_25_n_48 & {in2[1]}));
 assign mul_22_25_n_290 = ~((mul_22_25_n_30 & {in1[17]}) | (mul_22_25_n_22 & {in2[18]}));
 assign mul_22_25_n_289 = ~(({in2[29]} | mul_22_25_n_50) & ({in1[15]} | mul_22_25_n_53));
 assign mul_22_25_n_288 = ((mul_22_25_n_22 & ~{in1[18]}) | ({in1[17]} & {in1[18]}));
 assign mul_22_25_n_287 = ((mul_22_25_n_48 & ~{in1[8]}) | ({in1[7]} & {in1[8]}));
 assign mul_22_25_n_286 = ((mul_22_25_n_50 & ~{in1[16]}) | ({in1[15]} & {in1[16]}));
 assign mul_22_25_n_285 = ((mul_22_25_n_47 & ~{in1[4]}) | ({in1[3]} & {in1[4]}));
 assign mul_22_25_n_284 = ((mul_22_25_n_20 & ~{in1[6]}) | ({in1[5]} & {in1[6]}));
 assign mul_22_25_n_283 = ((mul_22_25_n_46 & ~{in1[10]}) | ({in1[9]} & {in1[10]}));
 assign mul_22_25_n_282 = ((mul_22_25_n_21 & ~{in1[14]}) | ({in1[13]} & {in1[14]}));
 assign mul_22_25_n_281 = ((mul_22_25_n_44 & ~{in1[2]}) | ({in1[1]} & {in1[2]}));
 assign mul_22_25_n_280 = ((mul_22_25_n_49 & ~{in1[12]}) | ({in1[11]} & {in1[12]}));
 assign mul_22_25_n_248 = ~mul_22_25_n_247;
 assign mul_22_25_n_175 = ~mul_22_25_n_174;
 assign mul_22_25_n_171 = ~mul_22_25_n_170;
 assign mul_22_25_n_138 = ~mul_22_25_n_137;
 assign mul_22_25_n_129 = ~mul_22_25_n_128;
 assign mul_22_25_n_104 = ~((mul_22_25_n_23 & {in1[5]}) | (mul_22_25_n_20 & {in2[0]}));
 assign mul_22_25_n_103 = ~((mul_22_25_n_23 & {in1[11]}) | (mul_22_25_n_49 & {in2[0]}));
 assign mul_22_25_n_102 = ~((mul_22_25_n_23 & {in1[3]}) | (mul_22_25_n_47 & {in2[0]}));
 assign mul_22_25_n_101 = ~((mul_22_25_n_23 & {in1[9]}) | (mul_22_25_n_46 & {in2[0]}));
 assign mul_22_25_n_100 = ~((mul_22_25_n_23 & {in1[13]}) | (mul_22_25_n_21 & {in2[0]}));
 assign mul_22_25_n_98 = ~((mul_22_25_n_23 & {in1[15]}) | (mul_22_25_n_50 & {in2[0]}));
 assign mul_22_25_n_97 = ~((mul_22_25_n_23 & {in1[7]}) | (mul_22_25_n_48 & {in2[0]}));
 assign mul_22_25_n_96 = ~((mul_22_25_n_23 & {in1[19]}) | (mul_22_25_n_45 & {in2[0]}));
 assign mul_22_25_n_95 = ~((mul_22_25_n_23 & {in1[17]}) | (mul_22_25_n_22 & {in2[0]}));
 assign mul_22_25_n_94 = ~(({in2[0]} | mul_22_25_n_44) & ({in1[1]} | mul_22_25_n_23));
 assign mul_22_25_n_269 = ~(({in2[23]} | mul_22_25_n_44) & ({in1[1]} | mul_22_25_n_60));
 assign mul_22_25_n_268 = ~((mul_22_25_n_39 & {in1[17]}) | (mul_22_25_n_22 & {in2[28]}));
 assign mul_22_25_n_267 = ~((mul_22_25_n_55 & {in1[13]}) | (mul_22_25_n_21 & {in2[20]}));
 assign mul_22_25_n_266 = ~((mul_22_25_n_37 & {in1[19]}) | (mul_22_25_n_45 & {in2[10]}));
 assign mul_22_25_n_265 = ~((mul_22_25_n_40 & {in1[17]}) | (mul_22_25_n_22 & {in2[15]}));
 assign mul_22_25_n_264 = ~((mul_22_25_n_27 & {in1[3]}) | (mul_22_25_n_47 & {in2[16]}));
 assign mul_22_25_n_263 = ~((mul_22_25_n_31 & {in1[13]}) | (mul_22_25_n_21 & {in2[9]}));
 assign mul_22_25_n_262 = ~((mul_22_25_n_28 & {in1[13]}) | (mul_22_25_n_21 & {in2[25]}));
 assign mul_22_25_n_261 = ~(({in2[20]} | mul_22_25_n_47) & ({in1[3]} | mul_22_25_n_55));
 assign mul_22_25_n_260 = ~(({in2[24]} | mul_22_25_n_47) & ({in1[3]} | mul_22_25_n_59));
 assign mul_22_25_n_259 = ~((mul_22_25_n_28 & {in1[7]}) | (mul_22_25_n_48 & {in2[25]}));
 assign mul_22_25_n_258 = ~((mul_22_25_n_60 & {in1[17]}) | (mul_22_25_n_22 & {in2[23]}));
 assign mul_22_25_n_257 = ~((mul_22_25_n_31 & {in1[3]}) | (mul_22_25_n_47 & {in2[9]}));
 assign mul_22_25_n_256 = ~((mul_22_25_n_40 & {in1[3]}) | (mul_22_25_n_47 & {in2[15]}));
 assign mul_22_25_n_255 = ~((mul_22_25_n_26 & {in1[9]}) | (mul_22_25_n_46 & {in2[12]}));
 assign mul_22_25_n_254 = ~((mul_22_25_n_31 & {in1[7]}) | (mul_22_25_n_48 & {in2[9]}));
 assign mul_22_25_n_253 = ~((mul_22_25_n_41 & {in1[3]}) | (mul_22_25_n_47 & {in2[13]}));
 assign mul_22_25_n_252 = ~((mul_22_25_n_59 & {in1[5]}) | (mul_22_25_n_20 & {in2[24]}));
 assign mul_22_25_n_251 = ~((mul_22_25_n_60 & {in1[15]}) | (mul_22_25_n_50 & {in2[23]}));
 assign mul_22_25_n_250 = ~((mul_22_25_n_35 & {in1[5]}) | (mul_22_25_n_20 & {in2[7]}));
 assign mul_22_25_n_249 = ~((mul_22_25_n_40 & {in1[13]}) | (mul_22_25_n_21 & {in2[15]}));
 assign mul_22_25_n_247 = ~(({in2[29]} | mul_22_25_n_21) & ({in1[13]} | mul_22_25_n_53));
 assign mul_22_25_n_246 = ~((mul_22_25_n_25 & {in1[9]}) | (mul_22_25_n_46 & {in2[4]}));
 assign mul_22_25_n_245 = ~((mul_22_25_n_60 & {in1[13]}) | (mul_22_25_n_21 & {in2[23]}));
 assign mul_22_25_n_244 = ~((mul_22_25_n_58 & {in1[9]}) | (mul_22_25_n_46 & {in2[3]}));
 assign mul_22_25_n_243 = ~((mul_22_25_n_36 & {in1[3]}) | (mul_22_25_n_47 & {in2[14]}));
 assign mul_22_25_n_242 = ~((mul_22_25_n_33 & {in1[17]}) | (mul_22_25_n_22 & {in2[17]}));
 assign mul_22_25_n_241 = ~((mul_22_25_n_38 & {in1[9]}) | (mul_22_25_n_46 & {in2[1]}));
 assign mul_22_25_n_240 = ~((mul_22_25_n_30 & {in1[7]}) | (mul_22_25_n_48 & {in2[18]}));
 assign mul_22_25_n_239 = ~(({in2[27]} | mul_22_25_n_44) & ({in1[1]} | mul_22_25_n_57));
 assign mul_22_25_n_238 = ~((mul_22_25_n_61 & {in1[9]}) | (mul_22_25_n_46 & {in2[22]}));
 assign mul_22_25_n_237 = ~((mul_22_25_n_33 & {in1[3]}) | (mul_22_25_n_47 & {in2[17]}));
 assign mul_22_25_n_236 = ~((mul_22_25_n_53 & {in1[7]}) | (mul_22_25_n_48 & {in2[29]}));
 assign mul_22_25_n_235 = ~((mul_22_25_n_60 & {in1[9]}) | (mul_22_25_n_46 & {in2[23]}));
 assign mul_22_25_n_234 = ~(({in2[26]} | mul_22_25_n_44) & ({in1[1]} | mul_22_25_n_24));
 assign mul_22_25_n_233 = ~((mul_22_25_n_58 & {in1[11]}) | (mul_22_25_n_49 & {in2[3]}));
 assign mul_22_25_n_232 = ~(({in2[28]} | mul_22_25_n_47) & ({in1[3]} | mul_22_25_n_39));
 assign mul_22_25_n_231 = ~((mul_22_25_n_32 & {in1[11]}) | (mul_22_25_n_49 & {in2[8]}));
 assign mul_22_25_n_230 = ~((mul_22_25_n_31 & {in1[5]}) | (mul_22_25_n_20 & {in2[9]}));
 assign mul_22_25_n_229 = ~(({in2[28]} | mul_22_25_n_50) & ({in1[15]} | mul_22_25_n_39));
 assign mul_22_25_n_228 = ~((mul_22_25_n_41 & {in1[13]}) | (mul_22_25_n_21 & {in2[13]}));
 assign mul_22_25_n_227 = ~((mul_22_25_n_35 & {in1[13]}) | (mul_22_25_n_21 & {in2[7]}));
 assign mul_22_25_n_226 = ~((mul_22_25_n_36 & {in1[17]}) | (mul_22_25_n_22 & {in2[14]}));
 assign mul_22_25_n_225 = ~((mul_22_25_n_54 & {in1[5]}) | (mul_22_25_n_20 & {in2[21]}));
 assign mul_22_25_n_224 = ~((mul_22_25_n_57 & {in1[9]}) | (mul_22_25_n_46 & {in2[27]}));
 assign mul_22_25_n_223 = ~((mul_22_25_n_57 & {in1[5]}) | (mul_22_25_n_20 & {in2[27]}));
 assign mul_22_25_n_222 = ~((mul_22_25_n_39 & {in1[11]}) | (mul_22_25_n_49 & {in2[28]}));
 assign mul_22_25_n_221 = ~((mul_22_25_n_61 & {in1[13]}) | (mul_22_25_n_21 & {in2[22]}));
 assign mul_22_25_n_220 = ~((mul_22_25_n_29 & {in1[13]}) | (mul_22_25_n_21 & {in2[2]}));
 assign mul_22_25_n_219 = ~((mul_22_25_n_56 & {in1[5]}) | (mul_22_25_n_20 & {in2[5]}));
 assign mul_22_25_n_218 = ~((mul_22_25_n_54 & {in1[11]}) | (mul_22_25_n_49 & {in2[21]}));
 assign mul_22_25_n_217 = ~((mul_22_25_n_32 & {in1[13]}) | (mul_22_25_n_21 & {in2[8]}));
 assign mul_22_25_n_216 = ~((mul_22_25_n_58 & {in1[15]}) | (mul_22_25_n_50 & {in2[3]}));
 assign mul_22_25_n_215 = ~((mul_22_25_n_33 & {in1[5]}) | (mul_22_25_n_20 & {in2[17]}));
 assign mul_22_25_n_214 = ~((mul_22_25_n_38 & {in1[3]}) | (mul_22_25_n_47 & {in2[1]}));
 assign mul_22_25_n_213 = ~(({in2[21]} | mul_22_25_n_44) & ({in1[1]} | mul_22_25_n_54));
 assign mul_22_25_n_212 = ~((mul_22_25_n_28 & {in1[15]}) | (mul_22_25_n_50 & {in2[25]}));
 assign mul_22_25_n_211 = ~(({in2[26]} | mul_22_25_n_47) & ({in1[3]} | mul_22_25_n_24));
 assign mul_22_25_n_210 = ~((mul_22_25_n_63 & {in1[3]}) | (mul_22_25_n_47 & {in2[6]}));
 assign mul_22_25_n_209 = ~((mul_22_25_n_34 & {in1[7]}) | (mul_22_25_n_48 & {in2[19]}));
 assign mul_22_25_n_208 = ~(({in2[28]} | mul_22_25_n_44) & ({in1[1]} | mul_22_25_n_39));
 assign mul_22_25_n_207 = ~((mul_22_25_n_27 & {in1[17]}) | (mul_22_25_n_22 & {in2[16]}));
 assign mul_22_25_n_206 = ~((mul_22_25_n_57 & {in1[17]}) | (mul_22_25_n_22 & {in2[27]}));
 assign mul_22_25_n_205 = ~(({in2[23]} | mul_22_25_n_47) & ({in1[3]} | mul_22_25_n_60));
 assign mul_22_25_n_204 = ~((mul_22_25_n_56 & {in1[17]}) | (mul_22_25_n_22 & {in2[5]}));
 assign mul_22_25_n_203 = ~((mul_22_25_n_33 & {in1[19]}) | (mul_22_25_n_45 & {in2[17]}));
 assign mul_22_25_n_202 = ~((mul_22_25_n_53 & {in1[11]}) | (mul_22_25_n_49 & {in2[29]}));
 assign mul_22_25_n_201 = ~((mul_22_25_n_62 & {in1[11]}) | (mul_22_25_n_49 & {in2[11]}));
 assign mul_22_25_n_200 = ~((mul_22_25_n_59 & {in1[15]}) | (mul_22_25_n_50 & {in2[24]}));
 assign mul_22_25_n_199 = ~((mul_22_25_n_55 & {in1[19]}) | (mul_22_25_n_45 & {in2[20]}));
 assign mul_22_25_n_198 = ~((mul_22_25_n_38 & {in1[15]}) | (mul_22_25_n_50 & {in2[1]}));
 assign mul_22_25_n_197 = ~((mul_22_25_n_34 & {in1[17]}) | (mul_22_25_n_22 & {in2[19]}));
 assign mul_22_25_n_196 = ~((mul_22_25_n_58 & {in1[17]}) | (mul_22_25_n_22 & {in2[3]}));
 assign mul_22_25_n_195 = ~((mul_22_25_n_25 & {in1[19]}) | (mul_22_25_n_45 & {in2[4]}));
 assign mul_22_25_n_194 = ~(({in2[24]} | mul_22_25_n_44) & ({in1[1]} | mul_22_25_n_59));
 assign mul_22_25_n_193 = ~((mul_22_25_n_41 & {in1[11]}) | (mul_22_25_n_49 & {in2[13]}));
 assign mul_22_25_n_192 = ~((mul_22_25_n_56 & {in1[3]}) | (mul_22_25_n_47 & {in2[5]}));
 assign mul_22_25_n_191 = ~((mul_22_25_n_61 & {in1[19]}) | (mul_22_25_n_45 & {in2[22]}));
 assign mul_22_25_n_190 = ~((mul_22_25_n_28 & {in1[11]}) | (mul_22_25_n_49 & {in2[25]}));
 assign mul_22_25_n_189 = ~((mul_22_25_n_41 & {in1[9]}) | (mul_22_25_n_46 & {in2[13]}));
 assign mul_22_25_n_188 = ~((mul_22_25_n_34 & {in1[15]}) | (mul_22_25_n_50 & {in2[19]}));
 assign mul_22_25_n_187 = ~((mul_22_25_n_24 & {in1[19]}) | (mul_22_25_n_45 & {in2[26]}));
 assign mul_22_25_n_186 = ~((mul_22_25_n_56 & {in1[7]}) | (mul_22_25_n_48 & {in2[5]}));
 assign mul_22_25_n_185 = ~((mul_22_25_n_63 & {in1[19]}) | (mul_22_25_n_45 & {in2[6]}));
 assign mul_22_25_n_184 = ~((mul_22_25_n_31 & {in1[9]}) | (mul_22_25_n_46 & {in2[9]}));
 assign mul_22_25_n_183 = ~((mul_22_25_n_26 & {in1[13]}) | (mul_22_25_n_21 & {in2[12]}));
 assign mul_22_25_n_182 = ~((mul_22_25_n_32 & {in1[7]}) | (mul_22_25_n_48 & {in2[8]}));
 assign mul_22_25_n_181 = ~((mul_22_25_n_35 & {in1[11]}) | (mul_22_25_n_49 & {in2[7]}));
 assign mul_22_25_n_180 = ~((mul_22_25_n_62 & {in1[15]}) | (mul_22_25_n_50 & {in2[11]}));
 assign mul_22_25_n_179 = ~((mul_22_25_n_55 & {in1[7]}) | (mul_22_25_n_48 & {in2[20]}));
 assign mul_22_25_n_178 = ~((mul_22_25_n_62 & {in1[5]}) | (mul_22_25_n_20 & {in2[11]}));
 assign mul_22_25_n_177 = ~((mul_22_25_n_39 & {in1[19]}) | (mul_22_25_n_45 & {in2[28]}));
 assign mul_22_25_n_176 = ~((mul_22_25_n_33 & {in1[9]}) | (mul_22_25_n_46 & {in2[17]}));
 assign mul_22_25_n_174 = ~(({in2[18]} | mul_22_25_n_47) & ({in1[3]} | mul_22_25_n_30));
 assign mul_22_25_n_173 = ~((mul_22_25_n_26 & {in1[7]}) | (mul_22_25_n_48 & {in2[12]}));
 assign mul_22_25_n_172 = ~(({in2[14]} | mul_22_25_n_44) & ({in1[1]} | mul_22_25_n_36));
 assign mul_22_25_n_170 = ~((mul_22_25_n_57 & {in1[13]}) | (mul_22_25_n_21 & {in2[27]}));
 assign mul_22_25_n_169 = ~((mul_22_25_n_35 & {in1[15]}) | (mul_22_25_n_50 & {in2[7]}));
 assign mul_22_25_n_168 = ~((mul_22_25_n_63 & {in1[15]}) | (mul_22_25_n_50 & {in2[6]}));
 assign mul_22_25_n_167 = ~((mul_22_25_n_62 & {in1[1]}) | (mul_22_25_n_44 & {in2[11]}));
 assign mul_22_25_n_166 = ~((mul_22_25_n_58 & {in1[19]}) | (mul_22_25_n_45 & {in2[3]}));
 assign mul_22_25_n_165 = ~((mul_22_25_n_25 & {in1[3]}) | (mul_22_25_n_47 & {in2[4]}));
 assign mul_22_25_n_164 = ~((mul_22_25_n_38 & {in1[11]}) | (mul_22_25_n_49 & {in2[1]}));
 assign mul_22_25_n_163 = ~((mul_22_25_n_40 & {in1[19]}) | (mul_22_25_n_45 & {in2[15]}));
 assign mul_22_25_n_162 = ~((mul_22_25_n_57 & {in1[19]}) | (mul_22_25_n_45 & {in2[27]}));
 assign mul_22_25_n_161 = ~(({in2[22]} | mul_22_25_n_47) & ({in1[3]} | mul_22_25_n_61));
 assign mul_22_25_n_160 = ~((mul_22_25_n_61 & {in1[5]}) | (mul_22_25_n_20 & {in2[22]}));
 assign mul_22_25_n_159 = ~((mul_22_25_n_26 & {in1[11]}) | (mul_22_25_n_49 & {in2[12]}));
 assign mul_22_25_n_158 = ~((mul_22_25_n_34 & {in1[19]}) | (mul_22_25_n_45 & {in2[19]}));
 assign mul_22_25_n_157 = ~((mul_22_25_n_32 & {in1[17]}) | (mul_22_25_n_22 & {in2[8]}));
 assign mul_22_25_n_156 = ~((mul_22_25_n_27 & {in1[15]}) | (mul_22_25_n_50 & {in2[16]}));
 assign mul_22_25_n_155 = ~((mul_22_25_n_38 & {in1[19]}) | (mul_22_25_n_45 & {in2[1]}));
 assign mul_22_25_n_154 = ~(({in2[25]} | mul_22_25_n_47) & ({in1[3]} | mul_22_25_n_28));
 assign mul_22_25_n_153 = ~(({in2[16]} | mul_22_25_n_44) & ({in1[1]} | mul_22_25_n_27));
 assign mul_22_25_n_152 = ~((mul_22_25_n_25 & {in1[5]}) | (mul_22_25_n_20 & {in2[4]}));
 assign mul_22_25_n_151 = ~((mul_22_25_n_27 & {in1[19]}) | (mul_22_25_n_45 & {in2[16]}));
 assign mul_22_25_n_150 = ~((mul_22_25_n_35 & {in1[17]}) | (mul_22_25_n_22 & {in2[7]}));
 assign mul_22_25_n_149 = ~((mul_22_25_n_36 & {in1[13]}) | (mul_22_25_n_21 & {in2[14]}));
 assign mul_22_25_n_148 = ~((mul_22_25_n_30 & {in1[11]}) | (mul_22_25_n_49 & {in2[18]}));
 assign mul_22_25_n_147 = ~((mul_22_25_n_36 & {in1[7]}) | (mul_22_25_n_48 & {in2[14]}));
 assign mul_22_25_n_146 = ~((mul_22_25_n_25 & {in1[13]}) | (mul_22_25_n_21 & {in2[4]}));
 assign mul_22_25_n_145 = ~((mul_22_25_n_55 & {in1[5]}) | (mul_22_25_n_20 & {in2[20]}));
 assign mul_22_25_n_144 = ~(({in2[27]} | mul_22_25_n_47) & ({in1[3]} | mul_22_25_n_57));
 assign mul_22_25_n_143 = ~((mul_22_25_n_53 & {in1[5]}) | (mul_22_25_n_20 & {in2[29]}));
 assign mul_22_25_n_142 = ~((mul_22_25_n_39 & {in1[9]}) | (mul_22_25_n_46 & {in2[28]}));
 assign mul_22_25_n_141 = ~((mul_22_25_n_62 & {in1[13]}) | (mul_22_25_n_21 & {in2[11]}));
 assign mul_22_25_n_140 = ~(({in2[29]} | mul_22_25_n_44) & ({in1[1]} | mul_22_25_n_53));
 assign mul_22_25_n_139 = ~((mul_22_25_n_62 & {in1[7]}) | (mul_22_25_n_48 & {in2[11]}));
 assign mul_22_25_n_137 = ~(({in2[27]} | mul_22_25_n_50) & ({in1[15]} | mul_22_25_n_57));
 assign mul_22_25_n_136 = ~((mul_22_25_n_24 & {in1[17]}) | (mul_22_25_n_22 & {in2[26]}));
 assign mul_22_25_n_135 = ~((mul_22_25_n_30 & {in1[13]}) | (mul_22_25_n_21 & {in2[18]}));
 assign mul_22_25_n_134 = ~(({in2[25]} | mul_22_25_n_44) & ({in1[1]} | mul_22_25_n_28));
 assign mul_22_25_n_133 = ~((mul_22_25_n_63 & {in1[13]}) | (mul_22_25_n_21 & {in2[6]}));
 assign mul_22_25_n_132 = ~((mul_22_25_n_32 & {in1[1]}) | (mul_22_25_n_44 & {in2[8]}));
 assign mul_22_25_n_131 = ~((mul_22_25_n_31 & {in1[19]}) | (mul_22_25_n_45 & {in2[9]}));
 assign mul_22_25_n_130 = ~((mul_22_25_n_24 & {in1[5]}) | (mul_22_25_n_20 & {in2[26]}));
 assign mul_22_25_n_128 = ~((mul_22_25_n_26 & {in1[1]}) | (mul_22_25_n_44 & {in2[12]}));
 assign mul_22_25_n_127 = ~((mul_22_25_n_41 & {in1[5]}) | (mul_22_25_n_20 & {in2[13]}));
 assign mul_22_25_n_126 = ~((mul_22_25_n_29 & {in1[11]}) | (mul_22_25_n_49 & {in2[2]}));
 assign mul_22_25_n_125 = ~((mul_22_25_n_63 & {in1[11]}) | (mul_22_25_n_49 & {in2[6]}));
 assign mul_22_25_n_124 = ~((mul_22_25_n_55 & {in1[9]}) | (mul_22_25_n_46 & {in2[20]}));
 assign mul_22_25_n_123 = ~((mul_22_25_n_29 & {in1[15]}) | (mul_22_25_n_50 & {in2[2]}));
 assign mul_22_25_n_122 = ~((mul_22_25_n_34 & {in1[9]}) | (mul_22_25_n_46 & {in2[19]}));
 assign mul_22_25_n_121 = ~((mul_22_25_n_53 & {in1[19]}) | (mul_22_25_n_45 & {in2[29]}));
 assign mul_22_25_n_120 = ~((mul_22_25_n_58 & {in1[3]}) | (mul_22_25_n_47 & {in2[3]}));
 assign mul_22_25_n_119 = ~((mul_22_25_n_32 & {in1[15]}) | (mul_22_25_n_50 & {in2[8]}));
 assign mul_22_25_n_118 = ~(({in2[1]} | mul_22_25_n_44) & ({in1[1]} | mul_22_25_n_38));
 assign mul_22_25_n_117 = ~((mul_22_25_n_40 & {in1[7]}) | (mul_22_25_n_48 & {in2[15]}));
 assign mul_22_25_n_116 = ~((mul_22_25_n_55 & {in1[15]}) | (mul_22_25_n_50 & {in2[20]}));
 assign mul_22_25_n_115 = ~((mul_22_25_n_61 & {in1[15]}) | (mul_22_25_n_50 & {in2[22]}));
 assign mul_22_25_n_114 = ~((mul_22_25_n_54 & {in1[15]}) | (mul_22_25_n_50 & {in2[21]}));
 assign mul_22_25_n_113 = ~((mul_22_25_n_28 & {in1[19]}) | (mul_22_25_n_45 & {in2[25]}));
 assign mul_22_25_n_112 = ~((mul_22_25_n_55 & {in1[17]}) | (mul_22_25_n_22 & {in2[20]}));
 assign mul_22_25_n_111 = ~((mul_22_25_n_25 & {in1[15]}) | (mul_22_25_n_50 & {in2[4]}));
 assign mul_22_25_n_110 = ~((mul_22_25_n_59 & {in1[9]}) | (mul_22_25_n_46 & {in2[24]}));
 assign mul_22_25_n_109 = ~((mul_22_25_n_58 & {in1[5]}) | (mul_22_25_n_20 & {in2[3]}));
 assign mul_22_25_n_108 = ~(({in2[22]} | mul_22_25_n_44) & ({in1[1]} | mul_22_25_n_61));
 assign mul_22_25_n_107 = ~((mul_22_25_n_41 & {in1[7]}) | (mul_22_25_n_48 & {in2[13]}));
 assign mul_22_25_n_106 = ~((mul_22_25_n_37 & {in1[7]}) | (mul_22_25_n_48 & {in2[10]}));
 assign mul_22_25_n_105 = (({in1[20]} | mul_22_25_n_45) & ({in1[19]} | mul_22_25_n_51));
 assign mul_22_25_n_92 = ~(mul_22_25_n_51 & {in2[19]});
 assign mul_22_25_n_91 = ~(mul_22_25_n_51 & {in2[12]});
 assign mul_22_25_n_90 = ~(mul_22_25_n_51 & {in2[26]});
 assign mul_22_25_n_89 = ~(mul_22_25_n_51 & {in2[20]});
 assign mul_22_25_n_88 = ~(mul_22_25_n_51 & {in2[28]});
 assign mul_22_25_n_87 = ~(mul_22_25_n_51 & {in2[14]});
 assign mul_22_25_n_86 = ~(mul_22_25_n_51 & {in2[27]});
 assign mul_22_25_n_85 = ~(mul_22_25_n_51 & {in2[11]});
 assign mul_22_25_n_84 = ~(mul_22_25_n_51 & {in2[7]});
 assign mul_22_25_n_83 = ~(mul_22_25_n_51 & {in2[8]});
 assign mul_22_25_n_82 = ~(mul_22_25_n_51 & {in2[15]});
 assign mul_22_25_n_81 = ~(mul_22_25_n_51 & {in2[5]});
 assign mul_22_25_n_80 = ~(mul_22_25_n_51 & {in2[2]});
 assign mul_22_25_n_79 = ~(mul_22_25_n_51 & {in2[23]});
 assign asc001_0_ = ~(mul_22_25_n_52 | mul_22_25_n_23);
 assign mul_22_25_n_78 = ~(mul_22_25_n_51 & {in2[22]});
 assign mul_22_25_n_77 = ~(mul_22_25_n_51 & {in2[3]});
 assign mul_22_25_n_76 = ~(mul_22_25_n_51 & {in2[10]});
 assign mul_22_25_n_75 = ~(mul_22_25_n_51 & {in2[17]});
 assign mul_22_25_n_74 = ~({in2[29]} | mul_22_25_n_51);
 assign mul_22_25_n_73 = ~(mul_22_25_n_51 & {in2[16]});
 assign mul_22_25_n_72 = ~(mul_22_25_n_51 & {in2[1]});
 assign mul_22_25_n_71 = ~(mul_22_25_n_51 & {in2[9]});
 assign mul_22_25_n_70 = ~(mul_22_25_n_51 & {in2[6]});
 assign mul_22_25_n_69 = ~(mul_22_25_n_51 & {in2[18]});
 assign mul_22_25_n_68 = ~(mul_22_25_n_51 & {in2[4]});
 assign mul_22_25_n_67 = ~(mul_22_25_n_51 & {in2[21]});
 assign mul_22_25_n_66 = ~(mul_22_25_n_51 & {in2[24]});
 assign mul_22_25_n_65 = ~(mul_22_25_n_51 & {in2[13]});
 assign mul_22_25_n_64 = ~(mul_22_25_n_51 & {in2[25]});
 assign mul_22_25_n_63 = ~{in2[6]};
 assign mul_22_25_n_62 = ~{in2[11]};
 assign mul_22_25_n_61 = ~{in2[22]};
 assign mul_22_25_n_60 = ~{in2[23]};
 assign mul_22_25_n_59 = ~{in2[24]};
 assign mul_22_25_n_58 = ~{in2[3]};
 assign mul_22_25_n_57 = ~{in2[27]};
 assign mul_22_25_n_56 = ~{in2[5]};
 assign mul_22_25_n_55 = ~{in2[20]};
 assign mul_22_25_n_54 = ~{in2[21]};
 assign mul_22_25_n_53 = ~{in2[29]};
 assign mul_22_25_n_52 = ~{in1[0]};
 assign mul_22_25_n_51 = ~{in1[20]};
 assign mul_22_25_n_50 = ~{in1[15]};
 assign mul_22_25_n_49 = ~{in1[11]};
 assign mul_22_25_n_48 = ~{in1[7]};
 assign mul_22_25_n_47 = ~{in1[3]};
 assign mul_22_25_n_46 = ~{in1[9]};
 assign mul_22_25_n_45 = ~{in1[19]};
 assign mul_22_25_n_44 = ~{in1[1]};
 assign mul_22_25_n_43 = ~{in2[30]};
 assign mul_22_25_n_42 = ~{in2[31]};
 assign mul_22_25_n_41 = ~{in2[13]};
 assign mul_22_25_n_40 = ~{in2[15]};
 assign mul_22_25_n_39 = ~{in2[28]};
 assign mul_22_25_n_38 = ~{in2[1]};
 assign mul_22_25_n_37 = ~{in2[10]};
 assign mul_22_25_n_36 = ~{in2[14]};
 assign mul_22_25_n_35 = ~{in2[7]};
 assign mul_22_25_n_34 = ~{in2[19]};
 assign mul_22_25_n_33 = ~{in2[17]};
 assign mul_22_25_n_32 = ~{in2[8]};
 assign mul_22_25_n_31 = ~{in2[9]};
 assign mul_22_25_n_30 = ~{in2[18]};
 assign mul_22_25_n_29 = ~{in2[2]};
 assign mul_22_25_n_28 = ~{in2[25]};
 assign mul_22_25_n_27 = ~{in2[16]};
 assign mul_22_25_n_26 = ~{in2[12]};
 assign mul_22_25_n_25 = ~{in2[4]};
 assign mul_22_25_n_24 = ~{in2[26]};
 assign mul_22_25_n_23 = ~{in2[0]};
 assign mul_22_25_n_22 = ~{in1[17]};
 assign mul_22_25_n_21 = ~{in1[13]};
 assign mul_22_25_n_20 = ~{in1[5]};
 assign asc001_48_ = ~(mul_22_25_n_970 ^ mul_22_25_n_1232);
 assign asc001_18_ = (mul_22_25_n_1050 ^ mul_22_25_n_1143);
 assign mul_22_25_n_16 = (n_150 | mul_22_25_n_1778);
 assign mul_22_25_n_15 = (mul_22_25_n_1762 & mul_22_25_n_1797);
 assign mul_22_25_n_14 = (mul_22_25_n_1760 | mul_22_25_n_1795);
 assign mul_22_25_n_13 = (mul_22_25_n_1774 | mul_22_25_n_1809);
 assign mul_22_25_n_12 = (mul_22_25_n_1782 | mul_22_25_n_1817);
 assign mul_22_25_n_11 = (mul_22_25_n_1754 & mul_22_25_n_1789);
 assign asc001_10_ = ~(mul_22_25_n_974 ^ mul_22_25_n_982);
 assign mul_22_25_n_9 = (mul_22_25_n_1266 | mul_22_25_n_1269);
 assign mul_22_25_n_8 = (mul_22_25_n_1750 & mul_22_25_n_1272);
 assign mul_22_25_n_7 = (mul_22_25_n_521 & ~(mul_22_25_n_484 & mul_22_25_n_435));
 assign mul_22_25_n_6 = (mul_22_25_n_517 & ~(mul_22_25_n_492 & mul_22_25_n_424));
 assign mul_22_25_n_5 = ~(mul_22_25_n_286 | ~mul_22_25_n_417);
 assign mul_22_25_n_4 = ~(~mul_22_25_n_287 & mul_22_25_n_431);
 assign mul_22_25_n_3 = ~(mul_22_25_n_285 | ~mul_22_25_n_429);
 assign mul_22_25_n_2 = ~(~mul_22_25_n_283 & mul_22_25_n_418);
 assign mul_22_25_n_1 = (mul_22_25_n_452 & ~(mul_22_25_n_451 & mul_22_25_n_430));
 assign mul_22_25_n_0 = ~(mul_22_25_n_3 | (~mul_22_25_n_423 & mul_22_25_n_488));
 assign n_0 = ~clr;
 assign n_210 = ~({in1[20]} & (~{in2[0]} & ~{in1[19]}));
 assign mul_22_25_n_1274 = (mul_22_25_n_1284 ^ (mul_22_25_n_469 ^ mul_22_25_n_803));
endmodule


