`timescale 1ps / 1ps
module fft2_Mul_32Sx32S_50S_4(
          in2,
          in1,
          out1,
          clk,
          clr
);
   input [31:0] in2;
   input [31:0] in1;
   output [49:0] out1;
   input clk;
   input clr;
wire mul_22_25_n_0, mul_22_25_n_1, mul_22_25_n_2, mul_22_25_n_3, mul_22_25_n_4,
     mul_22_25_n_5, mul_22_25_n_6, mul_22_25_n_7, mul_22_25_n_9, mul_22_25_n_10,
     mul_22_25_n_11, mul_22_25_n_12, mul_22_25_n_13, mul_22_25_n_15,
     mul_22_25_n_17, mul_22_25_n_18, mul_22_25_n_19, mul_22_25_n_20,
     mul_22_25_n_21, mul_22_25_n_22, mul_22_25_n_23, mul_22_25_n_24,
     mul_22_25_n_25, mul_22_25_n_26, mul_22_25_n_27, mul_22_25_n_28,
     mul_22_25_n_29, mul_22_25_n_30, mul_22_25_n_31, mul_22_25_n_32,
     mul_22_25_n_33, mul_22_25_n_34, mul_22_25_n_35, mul_22_25_n_36,
     mul_22_25_n_37, mul_22_25_n_38, mul_22_25_n_39, mul_22_25_n_40,
     mul_22_25_n_41, mul_22_25_n_42, mul_22_25_n_43, mul_22_25_n_44,
     mul_22_25_n_45, mul_22_25_n_46, mul_22_25_n_47, mul_22_25_n_48,
     mul_22_25_n_49, mul_22_25_n_50, mul_22_25_n_51, mul_22_25_n_52,
     mul_22_25_n_53, mul_22_25_n_54, mul_22_25_n_55, mul_22_25_n_56,
     mul_22_25_n_57, mul_22_25_n_58, mul_22_25_n_59, mul_22_25_n_60,
     mul_22_25_n_61, mul_22_25_n_62, mul_22_25_n_63, mul_22_25_n_64,
     mul_22_25_n_65, mul_22_25_n_67, mul_22_25_n_68, mul_22_25_n_69,
     mul_22_25_n_70, mul_22_25_n_71, mul_22_25_n_72, mul_22_25_n_73,
     mul_22_25_n_74, mul_22_25_n_75, mul_22_25_n_77, mul_22_25_n_78,
     mul_22_25_n_79, mul_22_25_n_80, mul_22_25_n_81, mul_22_25_n_82,
     mul_22_25_n_83, mul_22_25_n_84, mul_22_25_n_85, mul_22_25_n_86,
     mul_22_25_n_87, mul_22_25_n_88, mul_22_25_n_89, mul_22_25_n_90,
     mul_22_25_n_91, mul_22_25_n_92, mul_22_25_n_93, mul_22_25_n_94,
     mul_22_25_n_95, mul_22_25_n_96, mul_22_25_n_97, mul_22_25_n_98,
     mul_22_25_n_99, mul_22_25_n_100, mul_22_25_n_101, mul_22_25_n_102,
     mul_22_25_n_103, mul_22_25_n_104, mul_22_25_n_105, mul_22_25_n_106,
     mul_22_25_n_107, mul_22_25_n_108, mul_22_25_n_109, mul_22_25_n_110,
     mul_22_25_n_111, mul_22_25_n_112, mul_22_25_n_113, mul_22_25_n_114,
     mul_22_25_n_115, mul_22_25_n_116, mul_22_25_n_117, mul_22_25_n_118,
     mul_22_25_n_119, mul_22_25_n_120, mul_22_25_n_121, mul_22_25_n_122,
     mul_22_25_n_123, mul_22_25_n_124, mul_22_25_n_125, mul_22_25_n_126,
     mul_22_25_n_127, mul_22_25_n_128, mul_22_25_n_129, mul_22_25_n_130,
     mul_22_25_n_131, mul_22_25_n_132, mul_22_25_n_133, mul_22_25_n_134,
     mul_22_25_n_135, mul_22_25_n_136, mul_22_25_n_137, mul_22_25_n_138,
     mul_22_25_n_139, mul_22_25_n_140, mul_22_25_n_141, mul_22_25_n_142,
     mul_22_25_n_143, mul_22_25_n_144, mul_22_25_n_145, mul_22_25_n_146,
     mul_22_25_n_147, mul_22_25_n_148, mul_22_25_n_149, mul_22_25_n_150,
     mul_22_25_n_151, mul_22_25_n_152, mul_22_25_n_153, mul_22_25_n_154,
     mul_22_25_n_155, mul_22_25_n_156, mul_22_25_n_157, mul_22_25_n_158,
     mul_22_25_n_159, mul_22_25_n_160, mul_22_25_n_161, mul_22_25_n_162,
     mul_22_25_n_163, mul_22_25_n_164, mul_22_25_n_165, mul_22_25_n_166,
     mul_22_25_n_167, mul_22_25_n_168, mul_22_25_n_169, mul_22_25_n_170,
     mul_22_25_n_171, mul_22_25_n_172, mul_22_25_n_173, mul_22_25_n_174,
     mul_22_25_n_175, mul_22_25_n_176, mul_22_25_n_177, mul_22_25_n_178,
     mul_22_25_n_179, mul_22_25_n_180, mul_22_25_n_181, mul_22_25_n_182,
     mul_22_25_n_183, mul_22_25_n_184, mul_22_25_n_185, mul_22_25_n_186,
     mul_22_25_n_187, mul_22_25_n_188, mul_22_25_n_189, mul_22_25_n_190,
     mul_22_25_n_191, mul_22_25_n_192, mul_22_25_n_193, mul_22_25_n_194,
     mul_22_25_n_195, mul_22_25_n_196, mul_22_25_n_197, mul_22_25_n_198,
     mul_22_25_n_199, mul_22_25_n_200, mul_22_25_n_201, mul_22_25_n_202,
     mul_22_25_n_203, mul_22_25_n_204, mul_22_25_n_205, mul_22_25_n_206,
     mul_22_25_n_207, mul_22_25_n_208, mul_22_25_n_209, mul_22_25_n_210,
     mul_22_25_n_211, mul_22_25_n_212, mul_22_25_n_213, mul_22_25_n_214,
     mul_22_25_n_215, mul_22_25_n_216, mul_22_25_n_217, mul_22_25_n_218,
     mul_22_25_n_219, mul_22_25_n_220, mul_22_25_n_221, mul_22_25_n_222,
     mul_22_25_n_223, mul_22_25_n_224, mul_22_25_n_225, mul_22_25_n_226,
     mul_22_25_n_227, mul_22_25_n_228, mul_22_25_n_229, mul_22_25_n_230,
     mul_22_25_n_231, mul_22_25_n_232, mul_22_25_n_233, mul_22_25_n_234,
     mul_22_25_n_235, mul_22_25_n_236, mul_22_25_n_237, mul_22_25_n_238,
     mul_22_25_n_239, mul_22_25_n_240, mul_22_25_n_241, mul_22_25_n_242,
     mul_22_25_n_243, mul_22_25_n_244, mul_22_25_n_245, mul_22_25_n_246,
     mul_22_25_n_247, mul_22_25_n_248, mul_22_25_n_249, mul_22_25_n_250,
     mul_22_25_n_251, mul_22_25_n_252, mul_22_25_n_253, mul_22_25_n_254,
     mul_22_25_n_255, mul_22_25_n_256, mul_22_25_n_257, mul_22_25_n_258,
     mul_22_25_n_259, mul_22_25_n_260, mul_22_25_n_261, mul_22_25_n_262,
     mul_22_25_n_263, mul_22_25_n_264, mul_22_25_n_265, mul_22_25_n_266,
     mul_22_25_n_267, mul_22_25_n_268, mul_22_25_n_269, mul_22_25_n_270,
     mul_22_25_n_271, mul_22_25_n_272, mul_22_25_n_273, mul_22_25_n_274,
     mul_22_25_n_275, mul_22_25_n_276, mul_22_25_n_277, mul_22_25_n_278,
     mul_22_25_n_279, mul_22_25_n_280, mul_22_25_n_281, mul_22_25_n_282,
     mul_22_25_n_283, mul_22_25_n_284, mul_22_25_n_285, mul_22_25_n_286,
     mul_22_25_n_287, mul_22_25_n_288, mul_22_25_n_289, mul_22_25_n_290,
     mul_22_25_n_291, mul_22_25_n_292, mul_22_25_n_293, mul_22_25_n_294,
     mul_22_25_n_295, mul_22_25_n_296, mul_22_25_n_297, mul_22_25_n_298,
     mul_22_25_n_299, mul_22_25_n_300, mul_22_25_n_301, mul_22_25_n_302,
     mul_22_25_n_303, mul_22_25_n_304, mul_22_25_n_305, mul_22_25_n_306,
     mul_22_25_n_307, mul_22_25_n_308, mul_22_25_n_309, mul_22_25_n_310,
     mul_22_25_n_311, mul_22_25_n_312, mul_22_25_n_313, mul_22_25_n_314,
     mul_22_25_n_315, mul_22_25_n_316, mul_22_25_n_317, mul_22_25_n_318,
     mul_22_25_n_319, mul_22_25_n_320, mul_22_25_n_321, mul_22_25_n_322,
     mul_22_25_n_323, mul_22_25_n_324, mul_22_25_n_325, mul_22_25_n_326,
     mul_22_25_n_327, mul_22_25_n_328, mul_22_25_n_329, mul_22_25_n_330,
     mul_22_25_n_331, mul_22_25_n_332, mul_22_25_n_333, mul_22_25_n_334,
     mul_22_25_n_335, mul_22_25_n_336, mul_22_25_n_337, mul_22_25_n_338,
     mul_22_25_n_339, mul_22_25_n_340, mul_22_25_n_341, mul_22_25_n_342,
     mul_22_25_n_343, mul_22_25_n_344, mul_22_25_n_345, mul_22_25_n_346,
     mul_22_25_n_347, mul_22_25_n_348, mul_22_25_n_349, mul_22_25_n_350,
     mul_22_25_n_351, mul_22_25_n_352, mul_22_25_n_353, mul_22_25_n_354,
     mul_22_25_n_355, mul_22_25_n_356, mul_22_25_n_357, mul_22_25_n_358,
     mul_22_25_n_359, mul_22_25_n_360, mul_22_25_n_361, mul_22_25_n_362,
     mul_22_25_n_363, mul_22_25_n_364, mul_22_25_n_365, mul_22_25_n_366,
     mul_22_25_n_367, mul_22_25_n_368, mul_22_25_n_369, mul_22_25_n_370,
     mul_22_25_n_371, mul_22_25_n_372, mul_22_25_n_373, mul_22_25_n_374,
     mul_22_25_n_375, mul_22_25_n_376, mul_22_25_n_377, mul_22_25_n_378,
     mul_22_25_n_379, mul_22_25_n_380, mul_22_25_n_381, mul_22_25_n_382,
     mul_22_25_n_383, mul_22_25_n_384, mul_22_25_n_385, mul_22_25_n_386,
     mul_22_25_n_387, mul_22_25_n_388, mul_22_25_n_389, mul_22_25_n_390,
     mul_22_25_n_391, mul_22_25_n_392, mul_22_25_n_393, mul_22_25_n_394,
     mul_22_25_n_395, mul_22_25_n_396, mul_22_25_n_397, mul_22_25_n_398,
     mul_22_25_n_399, mul_22_25_n_400, mul_22_25_n_401, mul_22_25_n_402,
     mul_22_25_n_403, mul_22_25_n_404, mul_22_25_n_405, mul_22_25_n_406,
     mul_22_25_n_407, mul_22_25_n_408, mul_22_25_n_409, mul_22_25_n_410,
     mul_22_25_n_411, mul_22_25_n_412, mul_22_25_n_413, mul_22_25_n_414,
     mul_22_25_n_415, mul_22_25_n_416, mul_22_25_n_417, mul_22_25_n_418,
     mul_22_25_n_419, mul_22_25_n_420, mul_22_25_n_421, mul_22_25_n_422,
     mul_22_25_n_423, mul_22_25_n_424, mul_22_25_n_425, mul_22_25_n_426,
     mul_22_25_n_427, mul_22_25_n_428, mul_22_25_n_429, mul_22_25_n_430,
     mul_22_25_n_431, mul_22_25_n_432, mul_22_25_n_433, mul_22_25_n_434,
     mul_22_25_n_435, mul_22_25_n_436, mul_22_25_n_437, mul_22_25_n_438,
     mul_22_25_n_439, mul_22_25_n_440, mul_22_25_n_441, mul_22_25_n_442,
     mul_22_25_n_443, mul_22_25_n_444, mul_22_25_n_445, mul_22_25_n_446,
     mul_22_25_n_447, mul_22_25_n_448, mul_22_25_n_449, mul_22_25_n_450,
     mul_22_25_n_451, mul_22_25_n_452, mul_22_25_n_453, mul_22_25_n_454,
     mul_22_25_n_455, mul_22_25_n_456, mul_22_25_n_457, mul_22_25_n_458,
     mul_22_25_n_459, mul_22_25_n_460, mul_22_25_n_461, mul_22_25_n_462,
     mul_22_25_n_463, mul_22_25_n_464, mul_22_25_n_465, mul_22_25_n_466,
     mul_22_25_n_467, mul_22_25_n_468, mul_22_25_n_469, mul_22_25_n_470,
     mul_22_25_n_471, mul_22_25_n_472, mul_22_25_n_473, mul_22_25_n_474,
     mul_22_25_n_475, mul_22_25_n_476, mul_22_25_n_477, mul_22_25_n_478,
     mul_22_25_n_479, mul_22_25_n_480, mul_22_25_n_481, mul_22_25_n_482,
     mul_22_25_n_483, mul_22_25_n_484, mul_22_25_n_485, mul_22_25_n_486,
     mul_22_25_n_487, mul_22_25_n_488, mul_22_25_n_489, mul_22_25_n_490,
     mul_22_25_n_491, mul_22_25_n_492, mul_22_25_n_493, mul_22_25_n_494,
     mul_22_25_n_495, mul_22_25_n_496, mul_22_25_n_497, mul_22_25_n_498,
     mul_22_25_n_499, mul_22_25_n_500, mul_22_25_n_501, mul_22_25_n_502,
     mul_22_25_n_503, mul_22_25_n_504, mul_22_25_n_505, mul_22_25_n_506,
     mul_22_25_n_507, mul_22_25_n_508, mul_22_25_n_509, mul_22_25_n_510,
     mul_22_25_n_511, mul_22_25_n_512, mul_22_25_n_513, mul_22_25_n_514,
     mul_22_25_n_515, mul_22_25_n_516, mul_22_25_n_517, mul_22_25_n_518,
     mul_22_25_n_519, mul_22_25_n_520, mul_22_25_n_521, mul_22_25_n_522,
     mul_22_25_n_523, mul_22_25_n_524, mul_22_25_n_525, mul_22_25_n_526,
     mul_22_25_n_527, mul_22_25_n_528, mul_22_25_n_529, mul_22_25_n_530,
     mul_22_25_n_531, mul_22_25_n_532, mul_22_25_n_533, mul_22_25_n_534,
     mul_22_25_n_535, mul_22_25_n_536, mul_22_25_n_537, mul_22_25_n_538,
     mul_22_25_n_539, mul_22_25_n_540, mul_22_25_n_541, mul_22_25_n_542,
     mul_22_25_n_543, mul_22_25_n_544, mul_22_25_n_545, mul_22_25_n_546,
     mul_22_25_n_547, mul_22_25_n_548, mul_22_25_n_549, mul_22_25_n_550,
     mul_22_25_n_551, mul_22_25_n_552, mul_22_25_n_553, mul_22_25_n_554,
     mul_22_25_n_555, mul_22_25_n_556, mul_22_25_n_557, mul_22_25_n_558,
     mul_22_25_n_559, mul_22_25_n_560, mul_22_25_n_561, mul_22_25_n_562,
     mul_22_25_n_563, mul_22_25_n_564, mul_22_25_n_565, mul_22_25_n_566,
     mul_22_25_n_567, mul_22_25_n_568, mul_22_25_n_569, mul_22_25_n_570,
     mul_22_25_n_571, mul_22_25_n_572, mul_22_25_n_573, mul_22_25_n_574,
     mul_22_25_n_575, mul_22_25_n_576, mul_22_25_n_577, mul_22_25_n_578,
     mul_22_25_n_579, mul_22_25_n_580, mul_22_25_n_581, mul_22_25_n_582,
     mul_22_25_n_583, mul_22_25_n_584, mul_22_25_n_585, mul_22_25_n_586,
     mul_22_25_n_587, mul_22_25_n_588, mul_22_25_n_589, mul_22_25_n_590,
     mul_22_25_n_591, mul_22_25_n_592, mul_22_25_n_593, mul_22_25_n_594,
     mul_22_25_n_595, mul_22_25_n_596, mul_22_25_n_597, mul_22_25_n_598,
     mul_22_25_n_599, mul_22_25_n_600, mul_22_25_n_601, mul_22_25_n_602,
     mul_22_25_n_603, mul_22_25_n_604, mul_22_25_n_605, mul_22_25_n_606,
     mul_22_25_n_607, mul_22_25_n_608, mul_22_25_n_609, mul_22_25_n_610,
     mul_22_25_n_611, mul_22_25_n_612, mul_22_25_n_613, mul_22_25_n_614,
     mul_22_25_n_615, mul_22_25_n_616, mul_22_25_n_617, mul_22_25_n_618,
     mul_22_25_n_619, mul_22_25_n_620, mul_22_25_n_621, mul_22_25_n_622,
     mul_22_25_n_623, mul_22_25_n_624, mul_22_25_n_625, mul_22_25_n_626,
     mul_22_25_n_627, mul_22_25_n_628, mul_22_25_n_629, mul_22_25_n_630,
     mul_22_25_n_631, mul_22_25_n_632, mul_22_25_n_633, mul_22_25_n_634,
     mul_22_25_n_635, mul_22_25_n_636, mul_22_25_n_637, mul_22_25_n_638,
     mul_22_25_n_639, mul_22_25_n_640, mul_22_25_n_641, mul_22_25_n_642,
     mul_22_25_n_643, mul_22_25_n_644, mul_22_25_n_645, mul_22_25_n_646,
     mul_22_25_n_647, mul_22_25_n_648, mul_22_25_n_649, mul_22_25_n_650,
     mul_22_25_n_651, mul_22_25_n_652, mul_22_25_n_653, mul_22_25_n_654,
     mul_22_25_n_655, mul_22_25_n_656, mul_22_25_n_657, mul_22_25_n_658,
     mul_22_25_n_659, mul_22_25_n_660, mul_22_25_n_661, mul_22_25_n_662,
     mul_22_25_n_663, mul_22_25_n_664, mul_22_25_n_665, mul_22_25_n_666,
     mul_22_25_n_667, mul_22_25_n_668, mul_22_25_n_669, mul_22_25_n_670,
     mul_22_25_n_671, mul_22_25_n_672, mul_22_25_n_673, mul_22_25_n_674,
     mul_22_25_n_675, mul_22_25_n_676, mul_22_25_n_677, mul_22_25_n_678,
     mul_22_25_n_679, mul_22_25_n_680, mul_22_25_n_681, mul_22_25_n_682,
     mul_22_25_n_683, mul_22_25_n_684, mul_22_25_n_685, mul_22_25_n_686,
     mul_22_25_n_687, mul_22_25_n_688, mul_22_25_n_689, mul_22_25_n_690,
     mul_22_25_n_691, mul_22_25_n_692, mul_22_25_n_693, mul_22_25_n_694,
     mul_22_25_n_695, mul_22_25_n_696, mul_22_25_n_697, mul_22_25_n_698,
     mul_22_25_n_699, mul_22_25_n_700, mul_22_25_n_701, mul_22_25_n_702,
     mul_22_25_n_703, mul_22_25_n_704, mul_22_25_n_705, mul_22_25_n_706,
     mul_22_25_n_707, mul_22_25_n_708, mul_22_25_n_709, mul_22_25_n_710,
     mul_22_25_n_711, mul_22_25_n_712, mul_22_25_n_713, mul_22_25_n_714,
     mul_22_25_n_715, mul_22_25_n_716, mul_22_25_n_717, mul_22_25_n_718,
     mul_22_25_n_719, mul_22_25_n_720, mul_22_25_n_721, mul_22_25_n_722,
     mul_22_25_n_723, mul_22_25_n_724, mul_22_25_n_725, mul_22_25_n_726,
     mul_22_25_n_727, mul_22_25_n_728, mul_22_25_n_729, mul_22_25_n_730,
     mul_22_25_n_731, mul_22_25_n_732, mul_22_25_n_733, mul_22_25_n_734,
     mul_22_25_n_735, mul_22_25_n_736, mul_22_25_n_737, mul_22_25_n_738,
     mul_22_25_n_739, mul_22_25_n_740, mul_22_25_n_741, mul_22_25_n_742,
     mul_22_25_n_743, mul_22_25_n_744, mul_22_25_n_745, mul_22_25_n_746,
     mul_22_25_n_747, mul_22_25_n_748, mul_22_25_n_749, mul_22_25_n_750,
     mul_22_25_n_751, mul_22_25_n_752, mul_22_25_n_753, mul_22_25_n_754,
     mul_22_25_n_755, mul_22_25_n_756, mul_22_25_n_757, mul_22_25_n_758,
     mul_22_25_n_759, mul_22_25_n_760, mul_22_25_n_761, mul_22_25_n_762,
     mul_22_25_n_763, mul_22_25_n_764, mul_22_25_n_765, mul_22_25_n_766,
     mul_22_25_n_767, mul_22_25_n_768, mul_22_25_n_769, mul_22_25_n_770,
     mul_22_25_n_771, mul_22_25_n_772, mul_22_25_n_773, mul_22_25_n_774,
     mul_22_25_n_775, mul_22_25_n_776, mul_22_25_n_777, mul_22_25_n_778,
     mul_22_25_n_779, mul_22_25_n_780, mul_22_25_n_781, mul_22_25_n_782,
     mul_22_25_n_783, mul_22_25_n_784, mul_22_25_n_785, mul_22_25_n_786,
     mul_22_25_n_787, mul_22_25_n_788, mul_22_25_n_789, mul_22_25_n_790,
     mul_22_25_n_791, mul_22_25_n_792, mul_22_25_n_793, mul_22_25_n_794,
     mul_22_25_n_795, mul_22_25_n_796, mul_22_25_n_797, mul_22_25_n_798,
     mul_22_25_n_799, mul_22_25_n_800, mul_22_25_n_801, mul_22_25_n_802,
     mul_22_25_n_803, mul_22_25_n_804, mul_22_25_n_805, mul_22_25_n_806,
     mul_22_25_n_807, mul_22_25_n_808, mul_22_25_n_809, mul_22_25_n_810,
     mul_22_25_n_811, mul_22_25_n_812, mul_22_25_n_813, mul_22_25_n_814,
     mul_22_25_n_815, mul_22_25_n_816, mul_22_25_n_817, mul_22_25_n_818,
     mul_22_25_n_819, mul_22_25_n_820, mul_22_25_n_821, mul_22_25_n_822,
     mul_22_25_n_823, mul_22_25_n_824, mul_22_25_n_825, mul_22_25_n_826,
     mul_22_25_n_827, mul_22_25_n_828, mul_22_25_n_829, mul_22_25_n_830,
     mul_22_25_n_831, mul_22_25_n_832, mul_22_25_n_833, mul_22_25_n_834,
     mul_22_25_n_835, mul_22_25_n_836, mul_22_25_n_837, mul_22_25_n_838,
     mul_22_25_n_839, mul_22_25_n_840, mul_22_25_n_841, mul_22_25_n_842,
     mul_22_25_n_843, mul_22_25_n_844, mul_22_25_n_845, mul_22_25_n_846,
     mul_22_25_n_847, mul_22_25_n_848, mul_22_25_n_849, mul_22_25_n_850,
     mul_22_25_n_851, mul_22_25_n_852, mul_22_25_n_853, mul_22_25_n_854,
     mul_22_25_n_855, mul_22_25_n_856, mul_22_25_n_857, mul_22_25_n_858,
     mul_22_25_n_859, mul_22_25_n_860, mul_22_25_n_861, mul_22_25_n_862,
     mul_22_25_n_863, mul_22_25_n_864, mul_22_25_n_865, mul_22_25_n_866,
     mul_22_25_n_867, mul_22_25_n_868, mul_22_25_n_869, mul_22_25_n_870,
     mul_22_25_n_871, mul_22_25_n_872, mul_22_25_n_873, mul_22_25_n_874,
     mul_22_25_n_875, mul_22_25_n_876, mul_22_25_n_877, mul_22_25_n_878,
     mul_22_25_n_879, mul_22_25_n_880, mul_22_25_n_881, mul_22_25_n_882,
     mul_22_25_n_883, mul_22_25_n_884, mul_22_25_n_885, mul_22_25_n_886,
     mul_22_25_n_887, mul_22_25_n_888, mul_22_25_n_889, mul_22_25_n_890,
     mul_22_25_n_891, mul_22_25_n_892, mul_22_25_n_893, mul_22_25_n_894,
     mul_22_25_n_895, mul_22_25_n_896, mul_22_25_n_897, mul_22_25_n_898,
     mul_22_25_n_899, mul_22_25_n_900, mul_22_25_n_901, mul_22_25_n_902,
     mul_22_25_n_903, mul_22_25_n_904, mul_22_25_n_905, mul_22_25_n_906,
     mul_22_25_n_907, mul_22_25_n_908, mul_22_25_n_909, mul_22_25_n_910,
     mul_22_25_n_911, mul_22_25_n_912, mul_22_25_n_913, mul_22_25_n_914,
     mul_22_25_n_915, mul_22_25_n_916, mul_22_25_n_917, mul_22_25_n_918,
     mul_22_25_n_919, mul_22_25_n_920, mul_22_25_n_921, mul_22_25_n_922,
     mul_22_25_n_923, mul_22_25_n_924, mul_22_25_n_925, mul_22_25_n_926,
     mul_22_25_n_927, mul_22_25_n_928, mul_22_25_n_929, mul_22_25_n_930,
     mul_22_25_n_931, mul_22_25_n_932, mul_22_25_n_933, mul_22_25_n_934,
     mul_22_25_n_935, mul_22_25_n_936, mul_22_25_n_937, mul_22_25_n_938,
     mul_22_25_n_939, mul_22_25_n_940, mul_22_25_n_941, mul_22_25_n_942,
     mul_22_25_n_943, mul_22_25_n_944, mul_22_25_n_945, mul_22_25_n_946,
     mul_22_25_n_947, mul_22_25_n_948, mul_22_25_n_949, mul_22_25_n_950,
     mul_22_25_n_951, mul_22_25_n_952, mul_22_25_n_953, mul_22_25_n_954,
     mul_22_25_n_955, mul_22_25_n_956, mul_22_25_n_957, mul_22_25_n_958,
     mul_22_25_n_959, mul_22_25_n_960, mul_22_25_n_961, mul_22_25_n_962,
     mul_22_25_n_963, mul_22_25_n_964, mul_22_25_n_965, mul_22_25_n_966,
     mul_22_25_n_967, mul_22_25_n_968, mul_22_25_n_969, mul_22_25_n_970,
     mul_22_25_n_971, mul_22_25_n_972, mul_22_25_n_973, mul_22_25_n_974,
     mul_22_25_n_975, mul_22_25_n_976, mul_22_25_n_977, mul_22_25_n_978,
     mul_22_25_n_979, mul_22_25_n_980, mul_22_25_n_981, mul_22_25_n_982,
     mul_22_25_n_983, mul_22_25_n_984, mul_22_25_n_985, mul_22_25_n_986,
     mul_22_25_n_987, mul_22_25_n_988, mul_22_25_n_989, mul_22_25_n_990,
     mul_22_25_n_991, mul_22_25_n_992, mul_22_25_n_993, mul_22_25_n_994,
     mul_22_25_n_995, mul_22_25_n_996, mul_22_25_n_997, mul_22_25_n_998,
     mul_22_25_n_999, mul_22_25_n_1000, mul_22_25_n_1001, mul_22_25_n_1002,
     mul_22_25_n_1003, mul_22_25_n_1004, mul_22_25_n_1005, mul_22_25_n_1006,
     mul_22_25_n_1007, mul_22_25_n_1008, mul_22_25_n_1009, mul_22_25_n_1010,
     mul_22_25_n_1011, mul_22_25_n_1012, mul_22_25_n_1013, mul_22_25_n_1014,
     mul_22_25_n_1015, mul_22_25_n_1016, mul_22_25_n_1017, mul_22_25_n_1018,
     mul_22_25_n_1019, mul_22_25_n_1020, mul_22_25_n_1021, mul_22_25_n_1022,
     mul_22_25_n_1023, mul_22_25_n_1024, mul_22_25_n_1025, mul_22_25_n_1026,
     mul_22_25_n_1027, mul_22_25_n_1028, mul_22_25_n_1029, mul_22_25_n_1030,
     mul_22_25_n_1031, mul_22_25_n_1032, mul_22_25_n_1033, mul_22_25_n_1034,
     mul_22_25_n_1035, mul_22_25_n_1036, mul_22_25_n_1037, mul_22_25_n_1038,
     mul_22_25_n_1039, mul_22_25_n_1040, mul_22_25_n_1041, mul_22_25_n_1042,
     mul_22_25_n_1043, mul_22_25_n_1044, mul_22_25_n_1045, mul_22_25_n_1046,
     mul_22_25_n_1047, mul_22_25_n_1048, mul_22_25_n_1049, mul_22_25_n_1050,
     mul_22_25_n_1051, mul_22_25_n_1052, mul_22_25_n_1053, mul_22_25_n_1054,
     mul_22_25_n_1055, mul_22_25_n_1056, mul_22_25_n_1057, mul_22_25_n_1058,
     mul_22_25_n_1059, mul_22_25_n_1060, mul_22_25_n_1061, mul_22_25_n_1062,
     mul_22_25_n_1063, mul_22_25_n_1064, mul_22_25_n_1065, mul_22_25_n_1066,
     mul_22_25_n_1067, mul_22_25_n_1068, mul_22_25_n_1069, mul_22_25_n_1070,
     mul_22_25_n_1071, mul_22_25_n_1072, mul_22_25_n_1073, mul_22_25_n_1074,
     mul_22_25_n_1075, mul_22_25_n_1076, mul_22_25_n_1077, mul_22_25_n_1078,
     mul_22_25_n_1079, mul_22_25_n_1080, mul_22_25_n_1081, mul_22_25_n_1082,
     mul_22_25_n_1083, mul_22_25_n_1084, mul_22_25_n_1085, mul_22_25_n_1086,
     mul_22_25_n_1087, mul_22_25_n_1088, mul_22_25_n_1089, mul_22_25_n_1090,
     mul_22_25_n_1091, mul_22_25_n_1092, mul_22_25_n_1093, mul_22_25_n_1094,
     mul_22_25_n_1095, mul_22_25_n_1096, mul_22_25_n_1097, mul_22_25_n_1098,
     mul_22_25_n_1099, mul_22_25_n_1100, mul_22_25_n_1101, mul_22_25_n_1102,
     mul_22_25_n_1103, mul_22_25_n_1104, mul_22_25_n_1105, mul_22_25_n_1106,
     mul_22_25_n_1107, mul_22_25_n_1108, mul_22_25_n_1109, mul_22_25_n_1110,
     mul_22_25_n_1111, mul_22_25_n_1112, mul_22_25_n_1113, mul_22_25_n_1114,
     mul_22_25_n_1115, mul_22_25_n_1116, mul_22_25_n_1117, mul_22_25_n_1118,
     mul_22_25_n_1119, mul_22_25_n_1120, mul_22_25_n_1121, mul_22_25_n_1122,
     mul_22_25_n_1123, mul_22_25_n_1124, mul_22_25_n_1125, mul_22_25_n_1126,
     mul_22_25_n_1127, mul_22_25_n_1128, mul_22_25_n_1129, mul_22_25_n_1130,
     mul_22_25_n_1131, mul_22_25_n_1132, mul_22_25_n_1133, mul_22_25_n_1134,
     mul_22_25_n_1135, mul_22_25_n_1136, mul_22_25_n_1137, mul_22_25_n_1138,
     mul_22_25_n_1139, mul_22_25_n_1140, mul_22_25_n_1141, mul_22_25_n_1142,
     mul_22_25_n_1143, mul_22_25_n_1144, mul_22_25_n_1145, mul_22_25_n_1146,
     mul_22_25_n_1147, mul_22_25_n_1148, mul_22_25_n_1149, mul_22_25_n_1150,
     mul_22_25_n_1152, mul_22_25_n_1153, mul_22_25_n_1154, mul_22_25_n_1155,
     mul_22_25_n_1156, mul_22_25_n_1157, mul_22_25_n_1158, mul_22_25_n_1159,
     mul_22_25_n_1160, mul_22_25_n_1161, mul_22_25_n_1162, mul_22_25_n_1163,
     mul_22_25_n_1164, mul_22_25_n_1165, mul_22_25_n_1166, mul_22_25_n_1167,
     mul_22_25_n_1168, mul_22_25_n_1169, mul_22_25_n_1170, mul_22_25_n_1171,
     mul_22_25_n_1172, mul_22_25_n_1173, mul_22_25_n_1174, mul_22_25_n_1175,
     mul_22_25_n_1176, mul_22_25_n_1177, mul_22_25_n_1178, mul_22_25_n_1180,
     mul_22_25_n_1181, mul_22_25_n_1182, mul_22_25_n_1183, mul_22_25_n_1184,
     mul_22_25_n_1186, mul_22_25_n_1187, mul_22_25_n_1188, mul_22_25_n_1189,
     mul_22_25_n_1190, mul_22_25_n_1191, mul_22_25_n_1193, mul_22_25_n_1194,
     mul_22_25_n_1195, mul_22_25_n_1196, mul_22_25_n_1197, mul_22_25_n_1199,
     mul_22_25_n_1200, mul_22_25_n_1201, mul_22_25_n_1202, mul_22_25_n_1203,
     mul_22_25_n_1204, mul_22_25_n_1205, mul_22_25_n_1206, mul_22_25_n_1207,
     mul_22_25_n_1208, mul_22_25_n_1209, mul_22_25_n_1211, mul_22_25_n_1212,
     mul_22_25_n_1214, mul_22_25_n_1215, mul_22_25_n_1216, mul_22_25_n_1217,
     mul_22_25_n_1219, mul_22_25_n_1220, mul_22_25_n_1221, mul_22_25_n_1222,
     mul_22_25_n_1223, mul_22_25_n_1224, mul_22_25_n_1225, mul_22_25_n_1226,
     mul_22_25_n_1227, mul_22_25_n_1228, mul_22_25_n_1229, mul_22_25_n_1230,
     mul_22_25_n_1231, mul_22_25_n_1232, mul_22_25_n_1233, mul_22_25_n_1234,
     mul_22_25_n_1236, mul_22_25_n_1237, mul_22_25_n_1238, mul_22_25_n_1239,
     mul_22_25_n_1240, mul_22_25_n_1241, mul_22_25_n_1242, mul_22_25_n_1243,
     mul_22_25_n_1244, mul_22_25_n_1245, mul_22_25_n_1246, mul_22_25_n_1247,
     mul_22_25_n_1250, mul_22_25_n_1251, mul_22_25_n_1252, mul_22_25_n_1253,
     mul_22_25_n_1254, mul_22_25_n_1255, mul_22_25_n_1256, mul_22_25_n_1257,
     mul_22_25_n_1258, mul_22_25_n_1259, mul_22_25_n_1260, mul_22_25_n_1261,
     mul_22_25_n_1262, mul_22_25_n_1263, mul_22_25_n_1264, mul_22_25_n_1265,
     mul_22_25_n_1266, mul_22_25_n_1267, mul_22_25_n_1268, mul_22_25_n_1269,
     mul_22_25_n_1270, mul_22_25_n_1271, mul_22_25_n_1273, mul_22_25_n_1274,
     mul_22_25_n_1275, mul_22_25_n_1276, mul_22_25_n_1277, mul_22_25_n_1278,
     mul_22_25_n_1280, mul_22_25_n_1281, mul_22_25_n_1282, mul_22_25_n_1283,
     mul_22_25_n_1284, mul_22_25_n_1285, mul_22_25_n_1286, mul_22_25_n_1287,
     mul_22_25_n_1288, mul_22_25_n_1289, mul_22_25_n_1290, mul_22_25_n_1291,
     mul_22_25_n_1292, mul_22_25_n_1293, mul_22_25_n_1294, mul_22_25_n_1295,
     mul_22_25_n_1297, mul_22_25_n_1298, mul_22_25_n_1299, mul_22_25_n_1300,
     mul_22_25_n_1301, mul_22_25_n_1302, mul_22_25_n_1303, mul_22_25_n_1304,
     mul_22_25_n_1305, mul_22_25_n_1306, mul_22_25_n_1307, mul_22_25_n_1308,
     mul_22_25_n_1309, mul_22_25_n_1310, mul_22_25_n_1311, mul_22_25_n_1312,
     mul_22_25_n_1313, mul_22_25_n_1314, mul_22_25_n_1315, mul_22_25_n_1316,
     mul_22_25_n_1317, mul_22_25_n_1318, mul_22_25_n_1319, mul_22_25_n_1320,
     mul_22_25_n_1321, mul_22_25_n_1322, mul_22_25_n_1323, mul_22_25_n_1324,
     mul_22_25_n_1325, mul_22_25_n_1326, mul_22_25_n_1327, mul_22_25_n_1329,
     mul_22_25_n_1330, mul_22_25_n_1331, mul_22_25_n_1332, mul_22_25_n_1333,
     mul_22_25_n_1334, mul_22_25_n_1335, mul_22_25_n_1336, mul_22_25_n_1337,
     mul_22_25_n_1338, mul_22_25_n_1339, mul_22_25_n_1340, mul_22_25_n_1341,
     mul_22_25_n_1342, mul_22_25_n_1343, mul_22_25_n_1344, mul_22_25_n_1345,
     mul_22_25_n_1346, mul_22_25_n_1347, mul_22_25_n_1348, mul_22_25_n_1349,
     mul_22_25_n_1350, mul_22_25_n_1351, mul_22_25_n_1352, mul_22_25_n_1353,
     mul_22_25_n_1354, mul_22_25_n_1357, mul_22_25_n_1358, mul_22_25_n_1359,
     mul_22_25_n_1360, mul_22_25_n_1361, mul_22_25_n_1362, mul_22_25_n_1363,
     mul_22_25_n_1364, mul_22_25_n_1365, mul_22_25_n_1366, mul_22_25_n_1367,
     mul_22_25_n_1369, mul_22_25_n_1370, mul_22_25_n_1371, mul_22_25_n_1372,
     mul_22_25_n_1373, mul_22_25_n_1375, mul_22_25_n_1376, mul_22_25_n_1377,
     mul_22_25_n_1378, mul_22_25_n_1379, mul_22_25_n_1380, mul_22_25_n_1381,
     mul_22_25_n_1382, mul_22_25_n_1383, mul_22_25_n_1384, mul_22_25_n_1385,
     mul_22_25_n_1386, mul_22_25_n_1387, mul_22_25_n_1388, mul_22_25_n_1389,
     mul_22_25_n_1390, mul_22_25_n_1391, mul_22_25_n_1392, mul_22_25_n_1393,
     mul_22_25_n_1394, mul_22_25_n_1395, mul_22_25_n_1396, mul_22_25_n_1397,
     mul_22_25_n_1398, mul_22_25_n_1399, mul_22_25_n_1400, mul_22_25_n_1401,
     mul_22_25_n_1402, mul_22_25_n_1403, mul_22_25_n_1404, mul_22_25_n_1405,
     mul_22_25_n_1406, mul_22_25_n_1407, mul_22_25_n_1408, mul_22_25_n_1409,
     mul_22_25_n_1410, mul_22_25_n_1411, mul_22_25_n_1414, mul_22_25_n_1415,
     mul_22_25_n_1416, mul_22_25_n_1417, mul_22_25_n_1418, mul_22_25_n_1419,
     mul_22_25_n_1420, mul_22_25_n_1421, mul_22_25_n_1422, mul_22_25_n_1423,
     mul_22_25_n_1424, mul_22_25_n_1425, mul_22_25_n_1426, mul_22_25_n_1427,
     mul_22_25_n_1428, mul_22_25_n_1429, mul_22_25_n_1430, mul_22_25_n_1431,
     mul_22_25_n_1432, mul_22_25_n_1433, mul_22_25_n_1434, mul_22_25_n_1435,
     mul_22_25_n_1436, mul_22_25_n_1437, mul_22_25_n_1438, mul_22_25_n_1442,
     mul_22_25_n_1443, mul_22_25_n_1444, mul_22_25_n_1445, mul_22_25_n_1446,
     mul_22_25_n_1447, mul_22_25_n_1448, mul_22_25_n_1449, mul_22_25_n_1450,
     mul_22_25_n_1451, mul_22_25_n_1452, mul_22_25_n_1453, mul_22_25_n_1454,
     mul_22_25_n_1455, mul_22_25_n_1456, mul_22_25_n_1457, mul_22_25_n_1458,
     mul_22_25_n_1459, mul_22_25_n_1460, mul_22_25_n_1461, mul_22_25_n_1462,
     mul_22_25_n_1463, mul_22_25_n_1467, mul_22_25_n_1468, mul_22_25_n_1469,
     mul_22_25_n_1470, mul_22_25_n_1471, mul_22_25_n_1472, mul_22_25_n_1473,
     mul_22_25_n_1475, mul_22_25_n_1476, mul_22_25_n_1477, mul_22_25_n_1479,
     mul_22_25_n_1480, mul_22_25_n_1481, mul_22_25_n_1482, mul_22_25_n_1483,
     mul_22_25_n_1487, mul_22_25_n_1488, mul_22_25_n_1489, mul_22_25_n_1491,
     mul_22_25_n_1492, mul_22_25_n_1493, mul_22_25_n_1494, mul_22_25_n_1498,
     mul_22_25_n_1500, mul_22_25_n_1504, mul_22_25_n_1505, mul_22_25_n_1506,
     mul_22_25_n_1511, mul_22_25_n_1514, mul_22_25_n_1515, mul_22_25_n_1516,
     mul_22_25_n_1517, mul_22_25_n_1518, mul_22_25_n_1519, mul_22_25_n_1520,
     mul_22_25_n_1521, mul_22_25_n_1522, mul_22_25_n_1523, mul_22_25_n_1524,
     mul_22_25_n_1525, mul_22_25_n_1526, mul_22_25_n_1527, mul_22_25_n_1528,
     mul_22_25_n_1529, mul_22_25_n_1530, mul_22_25_n_1531, mul_22_25_n_1532,
     mul_22_25_n_1533, mul_22_25_n_1534, mul_22_25_n_1535, mul_22_25_n_1536,
     mul_22_25_n_1537, mul_22_25_n_1538, mul_22_25_n_1539, mul_22_25_n_1540,
     mul_22_25_n_1541, mul_22_25_n_1542, mul_22_25_n_1543, mul_22_25_n_1544,
     mul_22_25_n_1545, mul_22_25_n_1546, mul_22_25_n_1547, mul_22_25_n_1548,
     mul_22_25_n_1549, mul_22_25_n_1550, mul_22_25_n_1551, mul_22_25_n_1552,
     mul_22_25_n_1553, mul_22_25_n_1554, mul_22_25_n_1555, mul_22_25_n_1556,
     mul_22_25_n_1557, mul_22_25_n_1558, mul_22_25_n_1559, mul_22_25_n_1560,
     mul_22_25_n_1561, mul_22_25_n_1562, mul_22_25_n_1563, mul_22_25_n_1564,
     mul_22_25_n_1565, mul_22_25_n_1566, mul_22_25_n_1567, mul_22_25_n_1568,
     mul_22_25_n_1569, mul_22_25_n_1570, mul_22_25_n_1571, mul_22_25_n_1572,
     mul_22_25_n_1573, mul_22_25_n_1574, mul_22_25_n_1575, mul_22_25_n_1576,
     mul_22_25_n_1577, mul_22_25_n_1578, mul_22_25_n_1579, mul_22_25_n_1580,
     mul_22_25_n_1581, mul_22_25_n_1582, mul_22_25_n_1583, mul_22_25_n_1584,
     mul_22_25_n_1585, mul_22_25_n_1586, mul_22_25_n_1587, mul_22_25_n_1588,
     mul_22_25_n_1589, mul_22_25_n_1590, mul_22_25_n_1591, mul_22_25_n_1592,
     mul_22_25_n_1593, mul_22_25_n_1594, mul_22_25_n_1595, mul_22_25_n_1596,
     mul_22_25_n_1597, mul_22_25_n_1598, mul_22_25_n_1599, mul_22_25_n_1600,
     mul_22_25_n_1601, mul_22_25_n_1602, mul_22_25_n_1603, mul_22_25_n_1604,
     mul_22_25_n_1605, mul_22_25_n_1606, mul_22_25_n_1607, mul_22_25_n_1608,
     mul_22_25_n_1609, mul_22_25_n_1610, mul_22_25_n_1611, mul_22_25_n_1612,
     mul_22_25_n_1613, mul_22_25_n_1614, mul_22_25_n_1615, mul_22_25_n_1616,
     mul_22_25_n_1617, mul_22_25_n_1618, mul_22_25_n_1619, mul_22_25_n_1620,
     mul_22_25_n_1621, mul_22_25_n_1622, mul_22_25_n_1623, mul_22_25_n_1624,
     mul_22_25_n_1625, mul_22_25_n_1626, mul_22_25_n_1627, mul_22_25_n_1628,
     mul_22_25_n_1629, mul_22_25_n_1630, mul_22_25_n_1631, mul_22_25_n_1632,
     mul_22_25_n_1633, mul_22_25_n_1634, mul_22_25_n_1635, mul_22_25_n_1636,
     mul_22_25_n_1637, mul_22_25_n_1638, mul_22_25_n_1639, mul_22_25_n_1640,
     mul_22_25_n_1641, mul_22_25_n_1642, mul_22_25_n_1643, mul_22_25_n_1644,
     mul_22_25_n_1645, mul_22_25_n_1646, mul_22_25_n_1647, mul_22_25_n_1648,
     mul_22_25_n_1649, mul_22_25_n_1650, mul_22_25_n_1651, mul_22_25_n_1652,
     mul_22_25_n_1653, mul_22_25_n_1654, mul_22_25_n_1655, mul_22_25_n_1656,
     mul_22_25_n_1657, mul_22_25_n_1658, mul_22_25_n_1659, mul_22_25_n_1660,
     mul_22_25_n_1661, mul_22_25_n_1662, mul_22_25_n_1663, mul_22_25_n_1664,
     mul_22_25_n_1665, mul_22_25_n_1666, mul_22_25_n_1667, mul_22_25_n_1668,
     mul_22_25_n_1669, mul_22_25_n_1670, mul_22_25_n_1671, mul_22_25_n_1672,
     mul_22_25_n_1673, mul_22_25_n_1674, mul_22_25_n_1675, mul_22_25_n_1676,
     mul_22_25_n_1677, mul_22_25_n_1678, mul_22_25_n_1679, mul_22_25_n_1680,
     mul_22_25_n_1681, mul_22_25_n_1682, mul_22_25_n_1683, mul_22_25_n_1684,
     mul_22_25_n_1685, mul_22_25_n_1686, mul_22_25_n_1687, mul_22_25_n_1688,
     mul_22_25_n_1689, mul_22_25_n_1690, mul_22_25_n_1691, mul_22_25_n_1692,
     mul_22_25_n_1693, mul_22_25_n_1694, mul_22_25_n_1695, mul_22_25_n_1696,
     mul_22_25_n_1697, mul_22_25_n_1698, mul_22_25_n_1699, mul_22_25_n_1700,
     mul_22_25_n_1701, mul_22_25_n_1702, mul_22_25_n_1703, mul_22_25_n_1704,
     mul_22_25_n_1705, mul_22_25_n_1706, mul_22_25_n_1707, mul_22_25_n_1708,
     mul_22_25_n_1709, mul_22_25_n_1710, mul_22_25_n_1711, mul_22_25_n_1712,
     mul_22_25_n_1713, mul_22_25_n_1714, mul_22_25_n_1715, mul_22_25_n_1716,
     mul_22_25_n_1717, mul_22_25_n_1718, mul_22_25_n_1719, mul_22_25_n_1720,
     mul_22_25_n_1721, mul_22_25_n_1722, mul_22_25_n_1723, mul_22_25_n_1724,
     mul_22_25_n_1725, mul_22_25_n_1726, mul_22_25_n_1727, mul_22_25_n_1728,
     mul_22_25_n_1729, mul_22_25_n_1730, mul_22_25_n_1731, mul_22_25_n_1732,
     mul_22_25_n_1733, mul_22_25_n_1734, mul_22_25_n_1735, mul_22_25_n_1736,
     mul_22_25_n_1737, mul_22_25_n_1738, mul_22_25_n_1739, mul_22_25_n_1740,
     mul_22_25_n_1741, mul_22_25_n_1742, mul_22_25_n_1743, mul_22_25_n_1744,
     mul_22_25_n_1745, mul_22_25_n_1746, mul_22_25_n_1747, mul_22_25_n_1748,
     mul_22_25_n_1749, mul_22_25_n_1750, mul_22_25_n_1751, mul_22_25_n_1752,
     mul_22_25_n_1753, mul_22_25_n_1754, mul_22_25_n_1755, mul_22_25_n_1756,
     mul_22_25_n_1757, mul_22_25_n_1758, mul_22_25_n_1759, mul_22_25_n_1760,
     mul_22_25_n_1761, mul_22_25_n_1762, mul_22_25_n_1763, mul_22_25_n_1764,
     mul_22_25_n_1765, mul_22_25_n_1766, mul_22_25_n_1767, mul_22_25_n_1768,
     mul_22_25_n_1769, mul_22_25_n_1770, mul_22_25_n_1771, mul_22_25_n_1772,
     mul_22_25_n_1773, mul_22_25_n_1774, mul_22_25_n_1775, mul_22_25_n_1776,
     mul_22_25_n_1777, mul_22_25_n_1778, mul_22_25_n_1779, mul_22_25_n_1780,
     mul_22_25_n_1781, mul_22_25_n_1782, mul_22_25_n_1783, mul_22_25_n_1784,
     mul_22_25_n_1785, mul_22_25_n_1786, mul_22_25_n_1787, mul_22_25_n_1788,
     mul_22_25_n_1789, mul_22_25_n_1790, mul_22_25_n_1791, mul_22_25_n_1792,
     mul_22_25_n_1793, mul_22_25_n_1794, mul_22_25_n_1795, mul_22_25_n_1796,
     mul_22_25_n_1797, mul_22_25_n_1798, mul_22_25_n_1799, mul_22_25_n_1800,
     mul_22_25_n_1801, mul_22_25_n_1802, mul_22_25_n_1803, mul_22_25_n_1804,
     mul_22_25_n_1805, mul_22_25_n_1806, mul_22_25_n_1807, mul_22_25_n_1808,
     mul_22_25_n_1809, mul_22_25_n_1810, mul_22_25_n_1811, mul_22_25_n_1812,
     mul_22_25_n_1813, mul_22_25_n_1814, mul_22_25_n_1815, mul_22_25_n_1816,
     mul_22_25_n_1817, mul_22_25_n_1818, mul_22_25_n_1819, mul_22_25_n_1820,
     mul_22_25_n_1821, mul_22_25_n_1822, mul_22_25_n_1823, mul_22_25_n_1824,
     mul_22_25_n_1825, mul_22_25_n_1826, mul_22_25_n_1827, mul_22_25_n_1828,
     mul_22_25_n_1829, mul_22_25_n_1830, mul_22_25_n_1831, mul_22_25_n_1832,
     mul_22_25_n_1833, mul_22_25_n_1834, mul_22_25_n_1835, mul_22_25_n_1836,
     mul_22_25_n_1837, mul_22_25_n_1838, mul_22_25_n_1839, mul_22_25_n_1840,
     mul_22_25_n_1841, mul_22_25_n_1842, mul_22_25_n_1843, mul_22_25_n_1844,
     mul_22_25_n_1845, mul_22_25_n_1846, mul_22_25_n_1847, mul_22_25_n_1848,
     mul_22_25_n_1849, mul_22_25_n_1850, mul_22_25_n_1851, mul_22_25_n_1852,
     mul_22_25_n_1853, mul_22_25_n_1854, mul_22_25_n_1855, mul_22_25_n_1856,
     mul_22_25_n_1857, mul_22_25_n_1858, mul_22_25_n_1859, mul_22_25_n_1860,
     mul_22_25_n_1861, mul_22_25_n_1862, mul_22_25_n_1863, mul_22_25_n_1864,
     mul_22_25_n_1865, mul_22_25_n_1866, mul_22_25_n_1867, mul_22_25_n_1868,
     mul_22_25_n_1869, mul_22_25_n_1870, mul_22_25_n_1871, mul_22_25_n_1872,
     mul_22_25_n_1873, mul_22_25_n_1874, mul_22_25_n_1875, mul_22_25_n_1876,
     mul_22_25_n_1877, mul_22_25_n_1878, mul_22_25_n_1879, mul_22_25_n_1880,
     mul_22_25_n_1881, mul_22_25_n_1882, mul_22_25_n_1883, mul_22_25_n_1884,
     mul_22_25_n_1885, mul_22_25_n_1886, mul_22_25_n_1887, mul_22_25_n_1888,
     mul_22_25_n_1889, mul_22_25_n_1890, mul_22_25_n_1891, mul_22_25_n_1892,
     mul_22_25_n_1893, mul_22_25_n_1894, mul_22_25_n_1895, mul_22_25_n_1896,
     mul_22_25_n_1897, mul_22_25_n_1898, mul_22_25_n_1899, mul_22_25_n_1900,
     mul_22_25_n_1901, mul_22_25_n_1902, mul_22_25_n_1903, mul_22_25_n_1904,
     mul_22_25_n_1905, mul_22_25_n_1906, mul_22_25_n_1907, mul_22_25_n_1908,
     mul_22_25_n_1909, mul_22_25_n_1910, mul_22_25_n_1911, mul_22_25_n_1912,
     mul_22_25_n_1913, mul_22_25_n_1914, mul_22_25_n_1915, mul_22_25_n_1916,
     mul_22_25_n_1917, mul_22_25_n_1918, mul_22_25_n_1919, mul_22_25_n_1920,
     mul_22_25_n_1921, mul_22_25_n_1922, mul_22_25_n_1923, mul_22_25_n_1924,
     mul_22_25_n_1925, mul_22_25_n_1926, mul_22_25_n_1927, mul_22_25_n_1928,
     mul_22_25_n_1929, mul_22_25_n_1930, mul_22_25_n_1931, mul_22_25_n_1932,
     mul_22_25_n_1933, mul_22_25_n_1934, mul_22_25_n_1935, mul_22_25_n_1936,
     mul_22_25_n_1937, mul_22_25_n_1938, mul_22_25_n_1939, mul_22_25_n_1940,
     mul_22_25_n_1941, mul_22_25_n_1942, mul_22_25_n_1943, mul_22_25_n_1944,
     mul_22_25_n_1945, mul_22_25_n_1946, mul_22_25_n_1947, mul_22_25_n_1948,
     mul_22_25_n_1949, mul_22_25_n_1950, mul_22_25_n_1951, mul_22_25_n_1952,
     mul_22_25_n_1953, mul_22_25_n_1954, mul_22_25_n_1955, mul_22_25_n_1956,
     mul_22_25_n_1957, mul_22_25_n_1958, mul_22_25_n_1959, mul_22_25_n_1960,
     mul_22_25_n_1961, mul_22_25_n_1962, mul_22_25_n_1963, mul_22_25_n_1964,
     mul_22_25_n_1965, mul_22_25_n_1966, mul_22_25_n_1967, mul_22_25_n_1968,
     mul_22_25_n_1969, mul_22_25_n_1970, mul_22_25_n_1971, mul_22_25_n_1972,
     mul_22_25_n_1973, mul_22_25_n_1974, mul_22_25_n_1975, mul_22_25_n_1976,
     mul_22_25_n_1977, mul_22_25_n_1978, mul_22_25_n_1979, mul_22_25_n_1980,
     mul_22_25_n_1981, mul_22_25_n_1982, mul_22_25_n_1983, mul_22_25_n_1984,
     mul_22_25_n_1985, mul_22_25_n_1986, mul_22_25_n_1987, mul_22_25_n_1988,
     mul_22_25_n_1989, mul_22_25_n_1990, mul_22_25_n_1991, mul_22_25_n_1992,
     mul_22_25_n_1993, mul_22_25_n_1994, mul_22_25_n_1995, mul_22_25_n_1996,
     mul_22_25_n_1997, mul_22_25_n_1998, mul_22_25_n_1999, mul_22_25_n_2000,
     mul_22_25_n_2001, mul_22_25_n_2002, mul_22_25_n_2003, mul_22_25_n_2004,
     mul_22_25_n_2005, mul_22_25_n_2006, mul_22_25_n_2007, mul_22_25_n_2008,
     mul_22_25_n_2009, mul_22_25_n_2010, mul_22_25_n_2011, mul_22_25_n_2012,
     mul_22_25_n_2013, mul_22_25_n_2014, mul_22_25_n_2015, mul_22_25_n_2016,
     mul_22_25_n_2017, mul_22_25_n_2018, mul_22_25_n_2019, mul_22_25_n_2020,
     mul_22_25_n_2021, mul_22_25_n_2022, mul_22_25_n_2023, mul_22_25_n_2024,
     mul_22_25_n_2025, mul_22_25_n_2026, mul_22_25_n_2027, mul_22_25_n_2028,
     mul_22_25_n_2029, mul_22_25_n_2030, mul_22_25_n_2031, mul_22_25_n_2032,
     mul_22_25_n_2033, mul_22_25_n_2034, mul_22_25_n_2035, mul_22_25_n_2036,
     mul_22_25_n_2037, mul_22_25_n_2038, mul_22_25_n_2039, mul_22_25_n_2040,
     mul_22_25_n_2041, mul_22_25_n_2042, mul_22_25_n_2043, mul_22_25_n_2044,
     mul_22_25_n_2045, mul_22_25_n_2046, mul_22_25_n_2047, mul_22_25_n_2048,
     mul_22_25_n_2049, mul_22_25_n_2050, mul_22_25_n_2051, mul_22_25_n_2052,
     mul_22_25_n_2053, mul_22_25_n_2054, mul_22_25_n_2055, mul_22_25_n_2056,
     mul_22_25_n_2057, mul_22_25_n_2058, mul_22_25_n_2059, mul_22_25_n_2060,
     mul_22_25_n_2061, mul_22_25_n_2062, mul_22_25_n_2063, mul_22_25_n_2064,
     mul_22_25_n_2065, mul_22_25_n_2066, mul_22_25_n_2067, mul_22_25_n_2068,
     mul_22_25_n_2069, mul_22_25_n_2070, mul_22_25_n_2071, mul_22_25_n_2072,
     mul_22_25_n_2073, mul_22_25_n_2074, mul_22_25_n_2075, mul_22_25_n_2076,
     mul_22_25_n_2077, mul_22_25_n_2078, mul_22_25_n_2079, mul_22_25_n_2080,
     mul_22_25_n_2081, mul_22_25_n_2082, mul_22_25_n_2083, mul_22_25_n_2084,
     mul_22_25_n_2085, mul_22_25_n_2086, mul_22_25_n_2087, mul_22_25_n_2088,
     mul_22_25_n_2089, mul_22_25_n_2090, mul_22_25_n_2091, mul_22_25_n_2092,
     mul_22_25_n_2093, mul_22_25_n_2094, mul_22_25_n_2095, mul_22_25_n_2096,
     mul_22_25_n_2097, mul_22_25_n_2098, mul_22_25_n_2099, mul_22_25_n_2100,
     mul_22_25_n_2101, mul_22_25_n_2102, mul_22_25_n_2103, mul_22_25_n_2104,
     mul_22_25_n_2105, mul_22_25_n_2106, mul_22_25_n_2107, mul_22_25_n_2108,
     mul_22_25_n_2109, mul_22_25_n_2110, mul_22_25_n_2111, mul_22_25_n_2112,
     mul_22_25_n_2113, mul_22_25_n_2114, mul_22_25_n_2115, mul_22_25_n_2116,
     mul_22_25_n_2117, mul_22_25_n_2118, mul_22_25_n_2119, mul_22_25_n_2120,
     mul_22_25_n_2121, mul_22_25_n_2122, mul_22_25_n_2123, mul_22_25_n_2124,
     mul_22_25_n_2125, mul_22_25_n_2126, mul_22_25_n_2127, mul_22_25_n_2128,
     mul_22_25_n_2129, mul_22_25_n_2130, mul_22_25_n_2131, mul_22_25_n_2132,
     mul_22_25_n_2133, mul_22_25_n_2134, mul_22_25_n_2135, mul_22_25_n_2136,
     mul_22_25_n_2137, mul_22_25_n_2138, mul_22_25_n_2139, mul_22_25_n_2140,
     mul_22_25_n_2141, mul_22_25_n_2142, mul_22_25_n_2143, mul_22_25_n_2144,
     mul_22_25_n_2145, mul_22_25_n_2146, mul_22_25_n_2147, mul_22_25_n_2148,
     mul_22_25_n_2149, mul_22_25_n_2150, mul_22_25_n_2151, mul_22_25_n_2152,
     mul_22_25_n_2153, mul_22_25_n_2154, mul_22_25_n_2155, mul_22_25_n_2156,
     mul_22_25_n_2157, mul_22_25_n_2158, mul_22_25_n_2159, mul_22_25_n_2160,
     mul_22_25_n_2161, mul_22_25_n_2162, mul_22_25_n_2163, mul_22_25_n_2164,
     mul_22_25_n_2165, mul_22_25_n_2166, mul_22_25_n_2167, mul_22_25_n_2168,
     mul_22_25_n_2169, mul_22_25_n_2170, mul_22_25_n_2171, mul_22_25_n_2172,
     mul_22_25_n_2173, mul_22_25_n_2174, mul_22_25_n_2175, mul_22_25_n_2176,
     mul_22_25_n_2177, mul_22_25_n_2178, mul_22_25_n_2179, mul_22_25_n_2180,
     mul_22_25_n_2181, mul_22_25_n_2182, mul_22_25_n_2183, mul_22_25_n_2184,
     mul_22_25_n_2185, mul_22_25_n_2186, mul_22_25_n_2187, mul_22_25_n_2188,
     mul_22_25_n_2189, mul_22_25_n_2190, mul_22_25_n_2191, mul_22_25_n_2192,
     mul_22_25_n_2193, mul_22_25_n_2194, mul_22_25_n_2195, mul_22_25_n_2196,
     mul_22_25_n_2197, mul_22_25_n_2198, mul_22_25_n_2199, mul_22_25_n_2200,
     mul_22_25_n_2201, mul_22_25_n_2202, mul_22_25_n_2203, mul_22_25_n_2204,
     mul_22_25_n_2205, mul_22_25_n_2206, mul_22_25_n_2207, mul_22_25_n_2208,
     mul_22_25_n_2209, mul_22_25_n_2210, mul_22_25_n_2211, mul_22_25_n_2212,
     mul_22_25_n_2213, mul_22_25_n_2214, mul_22_25_n_2215, mul_22_25_n_2216,
     mul_22_25_n_2217, mul_22_25_n_2218, mul_22_25_n_2219, mul_22_25_n_2220,
     mul_22_25_n_2221, mul_22_25_n_2222, mul_22_25_n_2223, mul_22_25_n_2224,
     mul_22_25_n_2225, mul_22_25_n_2226, mul_22_25_n_2227, mul_22_25_n_2228,
     mul_22_25_n_2229, mul_22_25_n_2230, mul_22_25_n_2231, mul_22_25_n_2232,
     mul_22_25_n_2233, mul_22_25_n_2234, mul_22_25_n_2235, mul_22_25_n_2236,
     mul_22_25_n_2237, mul_22_25_n_2238, mul_22_25_n_2239, mul_22_25_n_2240,
     mul_22_25_n_2241, mul_22_25_n_2242, mul_22_25_n_2243, mul_22_25_n_2244,
     mul_22_25_n_2245, mul_22_25_n_2246, mul_22_25_n_2247, mul_22_25_n_2248,
     mul_22_25_n_2249, mul_22_25_n_2250, mul_22_25_n_2251, mul_22_25_n_2252,
     mul_22_25_n_2253, mul_22_25_n_2254, mul_22_25_n_2255, mul_22_25_n_2256,
     mul_22_25_n_2257, mul_22_25_n_2258, mul_22_25_n_2259, mul_22_25_n_2260,
     mul_22_25_n_2261, mul_22_25_n_2262, mul_22_25_n_2263, mul_22_25_n_2264,
     mul_22_25_n_2265, mul_22_25_n_2266, mul_22_25_n_2267, mul_22_25_n_2268,
     mul_22_25_n_2269, mul_22_25_n_2270, mul_22_25_n_2271, mul_22_25_n_2272,
     mul_22_25_n_2273, mul_22_25_n_2274, mul_22_25_n_2275, mul_22_25_n_2276,
     mul_22_25_n_2277, mul_22_25_n_2278, mul_22_25_n_2279, mul_22_25_n_2280,
     mul_22_25_n_2281, mul_22_25_n_2282, mul_22_25_n_2283, mul_22_25_n_2284,
     mul_22_25_n_2285, mul_22_25_n_2286, mul_22_25_n_2287, mul_22_25_n_2288,
     mul_22_25_n_2289, mul_22_25_n_2290, mul_22_25_n_2291, mul_22_25_n_2292,
     mul_22_25_n_2293, mul_22_25_n_2294, mul_22_25_n_2295, mul_22_25_n_2296,
     mul_22_25_n_2297, mul_22_25_n_2298, mul_22_25_n_2299, mul_22_25_n_2300,
     mul_22_25_n_2301, mul_22_25_n_2302, mul_22_25_n_2303, n_0, n_43, n_44, n_45,
     n_46, n_47, n_48, n_49, n_50, n_51, n_52, n_54, n_55, n_56, n_57, n_58,
     n_59, n_60, n_61, n_63, n_64, n_65, n_66, n_67, n_68, n_69, n_70, n_71,
     n_72, n_73, n_74, n_75, n_76, n_77, n_78, n_79, n_81, n_83, n_84, n_85,
     n_86, n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97,
     n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108,
     n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118, n_119,
     n_120, n_121, n_122, n_123, n_125, n_126, n_127, n_128, n_129, n_131, n_132,
     n_133, n_134, n_135, n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144,
     n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154, n_155,
     n_156, n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166,
     n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175, clk, clr, asc001_0_,
     asc001_1_, asc001_2_, asc001_3_, asc001_4_, asc001_5_, asc001_6_, asc001_7_,
     asc001_8_, asc001_9_, asc001_10_, asc001_11_, asc001_12_, asc001_13_,
     asc001_14_, asc001_15_, asc001_16_, asc001_17_, asc001_18_, asc001_19_,
     asc001_20_, asc001_21_, asc001_22_, asc001_23_, asc001_24_, asc001_25_,
     asc001_26_, asc001_27_, asc001_28_, asc001_29_, asc001_30_, asc001_31_,
     asc001_32_, asc001_33_, asc001_34_, asc001_35_, asc001_36_, asc001_37_,
     asc001_38_, asc001_39_, asc001_40_, asc001_41_, asc001_42_, asc001_43_,
     asc001_44_, asc001_45_, asc001_46_, asc001_47_, asc001_48_, asc001_49_;
assign {out1[49]} = asc001_49_;
assign {out1[48]} = asc001_48_;
assign {out1[47]} = asc001_47_;
assign {out1[46]} = asc001_46_;
assign {out1[45]} = asc001_45_;
assign {out1[44]} = asc001_44_;
assign {out1[43]} = asc001_43_;
assign {out1[42]} = asc001_42_;
assign {out1[41]} = asc001_41_;
assign {out1[40]} = asc001_40_;
assign {out1[39]} = asc001_39_;
assign {out1[38]} = asc001_38_;
assign {out1[37]} = asc001_37_;
assign {out1[36]} = asc001_36_;
assign {out1[35]} = asc001_35_;
assign {out1[34]} = asc001_34_;
assign {out1[33]} = asc001_33_;
assign {out1[32]} = asc001_32_;
assign {out1[31]} = asc001_31_;
assign {out1[30]} = asc001_30_;
assign {out1[29]} = asc001_29_;
assign {out1[28]} = asc001_28_;
assign {out1[27]} = asc001_27_;
assign {out1[26]} = asc001_26_;
assign {out1[25]} = asc001_25_;
assign {out1[24]} = asc001_24_;
assign {out1[23]} = asc001_23_;
assign {out1[22]} = asc001_22_;
assign {out1[21]} = asc001_21_;
assign {out1[20]} = asc001_20_;
assign {out1[19]} = asc001_19_;
assign {out1[18]} = asc001_18_;
assign {out1[17]} = asc001_17_;
assign {out1[16]} = asc001_16_;
assign {out1[15]} = asc001_15_;
assign {out1[14]} = asc001_14_;
assign {out1[13]} = asc001_13_;
assign {out1[12]} = asc001_12_;
assign {out1[11]} = asc001_11_;
assign {out1[10]} = asc001_10_;
assign {out1[9]} = asc001_9_;
 reg out1_41_L0_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) out1_41_L0_reg_IQ <= 1'B0;
     else begin
         out1_41_L0_reg_IQ <= asc001_8_;
     end
 assign {out1[8]} = out1_41_L0_reg_IQ;
 reg out1_42_L0_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) out1_42_L0_reg_IQ <= 1'B0;
     else begin
         out1_42_L0_reg_IQ <= asc001_7_;
     end
 assign {out1[7]} = out1_42_L0_reg_IQ;
 reg out1_43_L0_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) out1_43_L0_reg_IQ <= 1'B0;
     else begin
         out1_43_L0_reg_IQ <= asc001_6_;
     end
 assign {out1[6]} = out1_43_L0_reg_IQ;
 reg out1_44_L0_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) out1_44_L0_reg_IQ <= 1'B0;
     else begin
         out1_44_L0_reg_IQ <= asc001_5_;
     end
 assign {out1[5]} = out1_44_L0_reg_IQ;
 reg out1_45_L0_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) out1_45_L0_reg_IQ <= 1'B0;
     else begin
         out1_45_L0_reg_IQ <= asc001_4_;
     end
 assign {out1[4]} = out1_45_L0_reg_IQ;
 reg out1_46_L0_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) out1_46_L0_reg_IQ <= 1'B0;
     else begin
         out1_46_L0_reg_IQ <= asc001_3_;
     end
 assign {out1[3]} = out1_46_L0_reg_IQ;
 reg out1_47_L0_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) out1_47_L0_reg_IQ <= 1'B0;
     else begin
         out1_47_L0_reg_IQ <= asc001_2_;
     end
 assign {out1[2]} = out1_47_L0_reg_IQ;
 reg out1_48_L0_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) out1_48_L0_reg_IQ <= 1'B0;
     else begin
         out1_48_L0_reg_IQ <= asc001_1_;
     end
 assign {out1[1]} = out1_48_L0_reg_IQ;
 reg out1_49_L0_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) out1_49_L0_reg_IQ <= 1'B0;
     else begin
         out1_49_L0_reg_IQ <= asc001_0_;
     end
 assign {out1[0]} = out1_49_L0_reg_IQ;
 reg retime_s1_1_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_1_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_1_reg_reg_IQ <= mul_22_25_n_1685;
     end
 assign n_175 = retime_s1_1_reg_reg_IQ;
 reg retime_s1_2_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_2_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_2_reg_reg_IQ <= mul_22_25_n_1705;
     end
 assign n_174 = retime_s1_2_reg_reg_IQ;
 reg retime_s1_3_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_3_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_3_reg_reg_IQ <= mul_22_25_n_1708;
     end
 assign n_173 = retime_s1_3_reg_reg_IQ;
 reg retime_s1_4_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_4_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_4_reg_reg_IQ <= mul_22_25_n_1730;
     end
 assign n_172 = retime_s1_4_reg_reg_IQ;
 reg retime_s1_5_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_5_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_5_reg_reg_IQ <= mul_22_25_n_2056;
     end
 assign n_171 = retime_s1_5_reg_reg_IQ;
 reg retime_s1_6_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_6_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_6_reg_reg_IQ <= mul_22_25_n_2074;
     end
 assign n_170 = retime_s1_6_reg_reg_IQ;
 reg retime_s1_7_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_7_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_7_reg_reg_IQ <= mul_22_25_n_1774;
     end
 assign n_169 = retime_s1_7_reg_reg_IQ;
 reg retime_s1_8_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_8_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_8_reg_reg_IQ <= mul_22_25_n_1799;
     end
 assign n_168 = retime_s1_8_reg_reg_IQ;
 reg retime_s1_9_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_9_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_9_reg_reg_IQ <= mul_22_25_n_2018;
     end
 assign n_166 = retime_s1_9_reg_reg_IQ;
 reg retime_s1_10_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_10_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_10_reg_reg_IQ <= mul_22_25_n_1974;
     end
 assign n_165 = retime_s1_10_reg_reg_IQ;
 reg retime_s1_11_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_11_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_11_reg_reg_IQ <= mul_22_25_n_1995;
     end
 assign n_164 = retime_s1_11_reg_reg_IQ;
 reg retime_s1_12_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_12_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_12_reg_reg_IQ <= mul_22_25_n_1827;
     end
 assign n_163 = retime_s1_12_reg_reg_IQ;
 reg retime_s1_13_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_13_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_13_reg_reg_IQ <= mul_22_25_n_1853;
     end
 assign n_162 = retime_s1_13_reg_reg_IQ;
 reg retime_s1_14_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_14_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_14_reg_reg_IQ <= mul_22_25_n_2092;
     end
 assign n_161 = retime_s1_14_reg_reg_IQ;
 reg retime_s1_15_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_15_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_15_reg_reg_IQ <= mul_22_25_n_1905;
     end
 assign n_160 = retime_s1_15_reg_reg_IQ;
 reg retime_s1_16_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_16_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_16_reg_reg_IQ <= mul_22_25_n_1851;
     end
 assign n_159 = retime_s1_16_reg_reg_IQ;
 reg retime_s1_17_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_17_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_17_reg_reg_IQ <= mul_22_25_n_1877;
     end
 assign n_158 = retime_s1_17_reg_reg_IQ;
 reg retime_s1_18_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_18_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_18_reg_reg_IQ <= mul_22_25_n_2038;
     end
 assign n_157 = retime_s1_18_reg_reg_IQ;
 reg retime_s1_19_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_19_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_19_reg_reg_IQ <= mul_22_25_n_1610;
     end
 assign n_156 = retime_s1_19_reg_reg_IQ;
 reg retime_s1_20_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_20_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_20_reg_reg_IQ <= mul_22_25_n_1577;
     end
 assign n_155 = retime_s1_20_reg_reg_IQ;
 reg retime_s1_21_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_21_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_21_reg_reg_IQ <= mul_22_25_n_1593;
     end
 assign n_154 = retime_s1_21_reg_reg_IQ;
 reg retime_s1_22_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_22_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_22_reg_reg_IQ <= mul_22_25_n_2073;
     end
 assign n_153 = retime_s1_22_reg_reg_IQ;
 reg retime_s1_23_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_23_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_23_reg_reg_IQ <= mul_22_25_n_2091;
     end
 assign n_152 = retime_s1_23_reg_reg_IQ;
 reg retime_s1_24_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_24_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_24_reg_reg_IQ <= mul_22_25_n_2057;
     end
 assign n_151 = retime_s1_24_reg_reg_IQ;
 reg retime_s1_25_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_25_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_25_reg_reg_IQ <= mul_22_25_n_2075;
     end
 assign n_150 = retime_s1_25_reg_reg_IQ;
 reg retime_s1_26_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_26_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_26_reg_reg_IQ <= mul_22_25_n_1687;
     end
 assign n_149 = retime_s1_26_reg_reg_IQ;
 reg retime_s1_27_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_27_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_27_reg_reg_IQ <= mul_22_25_n_1707;
     end
 assign n_148 = retime_s1_27_reg_reg_IQ;
 reg retime_s1_28_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_28_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_28_reg_reg_IQ <= mul_22_25_n_1728;
     end
 assign n_147 = retime_s1_28_reg_reg_IQ;
 reg retime_s1_29_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_29_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_29_reg_reg_IQ <= mul_22_25_n_1751;
     end
 assign n_146 = retime_s1_29_reg_reg_IQ;
 reg retime_s1_30_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_30_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_30_reg_reg_IQ <= mul_22_25_n_2036;
     end
 assign n_145 = retime_s1_30_reg_reg_IQ;
 reg retime_s1_31_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_31_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_31_reg_reg_IQ <= mul_22_25_n_2055;
     end
 assign n_144 = retime_s1_31_reg_reg_IQ;
 reg retime_s1_32_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_32_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_32_reg_reg_IQ <= mul_22_25_n_1550;
     end
 assign n_143 = retime_s1_32_reg_reg_IQ;
 reg retime_s1_33_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_33_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_33_reg_reg_IQ <= mul_22_25_n_1564;
     end
 assign n_142 = retime_s1_33_reg_reg_IQ;
 reg retime_s1_34_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_34_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_34_reg_reg_IQ <= mul_22_25_n_1750;
     end
 assign n_141 = retime_s1_34_reg_reg_IQ;
 reg retime_s1_35_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_35_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_35_reg_reg_IQ <= mul_22_25_n_1775;
     end
 assign n_140 = retime_s1_35_reg_reg_IQ;
 reg retime_s1_36_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_36_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_36_reg_reg_IQ <= mul_22_25_n_2017;
     end
 assign n_139 = retime_s1_36_reg_reg_IQ;
 reg retime_s1_37_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_37_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_37_reg_reg_IQ <= mul_22_25_n_2037;
     end
 assign n_138 = retime_s1_37_reg_reg_IQ;
 reg retime_s1_38_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_38_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_38_reg_reg_IQ <= mul_22_25_n_2303;
     end
 assign n_137 = retime_s1_38_reg_reg_IQ;
 reg retime_s1_39_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_39_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_39_reg_reg_IQ <= mul_22_25_n_2270;
     end
 assign n_135 = retime_s1_39_reg_reg_IQ;
 reg retime_s1_40_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_40_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_40_reg_reg_IQ <= mul_22_25_n_1643;
     end
 assign n_134 = retime_s1_40_reg_reg_IQ;
 reg retime_s1_41_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_41_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_41_reg_reg_IQ <= mul_22_25_n_1663;
     end
 assign n_133 = retime_s1_41_reg_reg_IQ;
 reg retime_s1_42_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_42_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_42_reg_reg_IQ <= mul_22_25_n_1625;
     end
 assign n_132 = retime_s1_42_reg_reg_IQ;
 reg retime_s1_43_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_43_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_43_reg_reg_IQ <= mul_22_25_n_1644;
     end
 assign n_131 = retime_s1_43_reg_reg_IQ;
 reg retime_s1_44_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_44_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_44_reg_reg_IQ <= mul_22_25_n_1997;
     end
 assign n_129 = retime_s1_44_reg_reg_IQ;
 reg retime_s1_45_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_45_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_45_reg_reg_IQ <= mul_22_25_n_1951;
     end
 assign n_128 = retime_s1_45_reg_reg_IQ;
 reg retime_s1_46_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_46_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_46_reg_reg_IQ <= mul_22_25_n_1973;
     end
 assign n_127 = retime_s1_46_reg_reg_IQ;
 reg retime_s1_47_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_47_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_47_reg_reg_IQ <= mul_22_25_n_1927;
     end
 assign n_126 = retime_s1_47_reg_reg_IQ;
 reg retime_s1_48_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_48_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_48_reg_reg_IQ <= mul_22_25_n_1950;
     end
 assign n_125 = retime_s1_48_reg_reg_IQ;
 reg retime_s1_49_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_49_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_49_reg_reg_IQ <= mul_22_25_n_1232;
     end
 assign n_123 = retime_s1_49_reg_reg_IQ;
 reg retime_s1_50_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_50_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_50_reg_reg_IQ <= mul_22_25_n_1217;
     end
 assign n_122 = retime_s1_50_reg_reg_IQ;
 reg retime_s1_51_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_51_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_51_reg_reg_IQ <= mul_22_25_n_1930;
     end
 assign n_121 = retime_s1_51_reg_reg_IQ;
 reg retime_s1_52_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_52_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_52_reg_reg_IQ <= mul_22_25_n_1776;
     end
 assign n_120 = retime_s1_52_reg_reg_IQ;
 reg retime_s1_53_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_53_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_53_reg_reg_IQ <= mul_22_25_n_1802;
     end
 assign n_119 = retime_s1_53_reg_reg_IQ;
 reg retime_s1_54_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_54_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_54_reg_reg_IQ <= mul_22_25_n_1800;
     end
 assign n_118 = retime_s1_54_reg_reg_IQ;
 reg retime_s1_55_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_55_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_55_reg_reg_IQ <= mul_22_25_n_1825;
     end
 assign n_117 = retime_s1_55_reg_reg_IQ;
 reg retime_s1_56_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_56_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_56_reg_reg_IQ <= mul_22_25_n_1594;
     end
 assign n_116 = retime_s1_56_reg_reg_IQ;
 reg retime_s1_57_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_57_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_57_reg_reg_IQ <= mul_22_25_n_1563;
     end
 assign n_115 = retime_s1_57_reg_reg_IQ;
 reg retime_s1_58_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_58_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_58_reg_reg_IQ <= mul_22_25_n_1578;
     end
 assign n_114 = retime_s1_58_reg_reg_IQ;
 reg retime_s1_59_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_59_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_59_reg_reg_IQ <= mul_22_25_n_1579;
     end
 assign n_113 = retime_s1_59_reg_reg_IQ;
 reg retime_s1_60_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_60_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_60_reg_reg_IQ <= mul_22_25_n_1552;
     end
 assign n_112 = retime_s1_60_reg_reg_IQ;
 reg retime_s1_61_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_61_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_61_reg_reg_IQ <= mul_22_25_n_1565;
     end
 assign n_111 = retime_s1_61_reg_reg_IQ;
 reg retime_s1_62_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_62_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_62_reg_reg_IQ <= mul_22_25_n_1931;
     end
 assign n_110 = retime_s1_62_reg_reg_IQ;
 reg retime_s1_63_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_63_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_63_reg_reg_IQ <= mul_22_25_n_1664;
     end
 assign n_109 = retime_s1_63_reg_reg_IQ;
 reg retime_s1_64_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_64_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_64_reg_reg_IQ <= mul_22_25_n_1627;
     end
 assign n_108 = retime_s1_64_reg_reg_IQ;
 reg retime_s1_65_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_65_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_65_reg_reg_IQ <= mul_22_25_n_1645;
     end
 assign n_107 = retime_s1_65_reg_reg_IQ;
 reg retime_s1_66_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_66_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_66_reg_reg_IQ <= mul_22_25_n_1906;
     end
 assign n_106 = retime_s1_66_reg_reg_IQ;
 reg retime_s1_67_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_67_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_67_reg_reg_IQ <= mul_22_25_n_1706;
     end
 assign n_105 = retime_s1_67_reg_reg_IQ;
 reg retime_s1_68_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_68_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_68_reg_reg_IQ <= mul_22_25_n_1727;
     end
 assign n_104 = retime_s1_68_reg_reg_IQ;
 reg retime_s1_69_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_69_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_69_reg_reg_IQ <= mul_22_25_n_1753;
     end
 assign n_103 = retime_s1_69_reg_reg_IQ;
 reg retime_s1_70_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_70_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_70_reg_reg_IQ <= mul_22_25_n_1777;
     end
 assign n_102 = retime_s1_70_reg_reg_IQ;
 reg retime_s1_71_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_71_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_71_reg_reg_IQ <= mul_22_25_n_1540;
     end
 assign n_101 = retime_s1_71_reg_reg_IQ;
 reg retime_s1_72_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_72_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_72_reg_reg_IQ <= mul_22_25_n_1880;
     end
 assign n_100 = retime_s1_72_reg_reg_IQ;
 reg retime_s1_73_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_73_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_73_reg_reg_IQ <= mul_22_25_n_1826;
     end
 assign n_99 = retime_s1_73_reg_reg_IQ;
 reg retime_s1_74_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_74_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_74_reg_reg_IQ <= mul_22_25_n_1852;
     end
 assign n_98 = retime_s1_74_reg_reg_IQ;
 reg retime_s1_75_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_75_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_75_reg_reg_IQ <= mul_22_25_n_1975;
     end
 assign n_97 = retime_s1_75_reg_reg_IQ;
 reg retime_s1_76_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_76_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_76_reg_reg_IQ <= mul_22_25_n_2231;
     end
 assign n_96 = retime_s1_76_reg_reg_IQ;
 reg retime_s1_77_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_77_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_77_reg_reg_IQ <= mul_22_25_n_1258;
     end
 assign n_95 = retime_s1_77_reg_reg_IQ;
 reg retime_s1_78_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_78_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_78_reg_reg_IQ <= mul_22_25_n_2233;
     end
 assign n_94 = retime_s1_78_reg_reg_IQ;
 reg retime_s1_79_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_79_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_79_reg_reg_IQ <= mul_22_25_n_1268;
     end
 assign n_93 = retime_s1_79_reg_reg_IQ;
 reg retime_s1_80_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_80_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_80_reg_reg_IQ <= mul_22_25_n_2122;
     end
 assign n_92 = retime_s1_80_reg_reg_IQ;
 reg retime_s1_81_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_81_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_81_reg_reg_IQ <= mul_22_25_n_1233;
     end
 assign n_91 = retime_s1_81_reg_reg_IQ;
 reg retime_s1_82_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_82_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_82_reg_reg_IQ <= mul_22_25_n_1226;
     end
 assign n_90 = retime_s1_82_reg_reg_IQ;
 reg retime_s1_83_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_83_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_83_reg_reg_IQ <= mul_22_25_n_1225;
     end
 assign n_89 = retime_s1_83_reg_reg_IQ;
 reg retime_s1_84_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_84_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_84_reg_reg_IQ <= mul_22_25_n_1238;
     end
 assign n_88 = retime_s1_84_reg_reg_IQ;
 reg retime_s1_85_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_85_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_85_reg_reg_IQ <= mul_22_25_n_1224;
     end
 assign n_87 = retime_s1_85_reg_reg_IQ;
 reg retime_s1_86_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_86_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_86_reg_reg_IQ <= mul_22_25_n_2272;
     end
 assign n_86 = retime_s1_86_reg_reg_IQ;
 reg retime_s1_87_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_87_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_87_reg_reg_IQ <= mul_22_25_n_1237;
     end
 assign n_85 = retime_s1_87_reg_reg_IQ;
 reg retime_s1_88_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_88_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_88_reg_reg_IQ <= mul_22_25_n_1252;
     end
 assign n_84 = retime_s1_88_reg_reg_IQ;
 reg retime_s1_89_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_89_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_89_reg_reg_IQ <= mul_22_25_n_1250;
     end
 assign n_83 = retime_s1_89_reg_reg_IQ;
 reg retime_s1_90_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_90_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_90_reg_reg_IQ <= mul_22_25_n_1257;
     end
 assign n_81 = retime_s1_90_reg_reg_IQ;
 reg retime_s1_91_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_91_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_91_reg_reg_IQ <= mul_22_25_n_1592;
     end
 assign n_79 = retime_s1_91_reg_reg_IQ;
 reg retime_s1_92_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_92_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_92_reg_reg_IQ <= mul_22_25_n_1609;
     end
 assign n_78 = retime_s1_92_reg_reg_IQ;
 reg retime_s1_93_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_93_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_93_reg_reg_IQ <= mul_22_25_n_1879;
     end
 assign n_77 = retime_s1_93_reg_reg_IQ;
 reg retime_s1_94_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_94_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_94_reg_reg_IQ <= mul_22_25_n_1801;
     end
 assign n_76 = retime_s1_94_reg_reg_IQ;
 reg retime_s1_95_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_95_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_95_reg_reg_IQ <= mul_22_25_n_1828;
     end
 assign n_75 = retime_s1_95_reg_reg_IQ;
 reg retime_s1_96_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_96_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_96_reg_reg_IQ <= mul_22_25_n_1928;
     end
 assign n_74 = retime_s1_96_reg_reg_IQ;
 reg retime_s1_97_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_97_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_97_reg_reg_IQ <= mul_22_25_n_1952;
     end
 assign n_73 = retime_s1_97_reg_reg_IQ;
 reg retime_s1_98_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_98_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_98_reg_reg_IQ <= mul_22_25_n_1996;
     end
 assign n_72 = retime_s1_98_reg_reg_IQ;
 reg retime_s1_99_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_99_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_99_reg_reg_IQ <= mul_22_25_n_2016;
     end
 assign n_71 = retime_s1_99_reg_reg_IQ;
 reg retime_s1_100_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_100_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_100_reg_reg_IQ <= mul_22_25_n_1904;
     end
 assign n_70 = retime_s1_100_reg_reg_IQ;
 reg retime_s1_101_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_101_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_101_reg_reg_IQ <= mul_22_25_n_1929;
     end
 assign n_69 = retime_s1_101_reg_reg_IQ;
 reg retime_s1_102_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_102_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_102_reg_reg_IQ <= mul_22_25_n_1854;
     end
 assign n_68 = retime_s1_102_reg_reg_IQ;
 reg retime_s1_103_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_103_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_103_reg_reg_IQ <= mul_22_25_n_2107;
     end
 assign n_67 = retime_s1_103_reg_reg_IQ;
 reg retime_s1_104_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_104_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_104_reg_reg_IQ <= mul_22_25_n_2121;
     end
 assign n_66 = retime_s1_104_reg_reg_IQ;
 reg retime_s1_105_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_105_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_105_reg_reg_IQ <= mul_22_25_n_1227;
     end
 assign n_65 = retime_s1_105_reg_reg_IQ;
 reg retime_s1_106_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_106_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_106_reg_reg_IQ <= mul_22_25_n_1878;
     end
 assign n_64 = retime_s1_106_reg_reg_IQ;
 reg retime_s1_107_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_107_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_107_reg_reg_IQ <= mul_22_25_n_1903;
     end
 assign n_63 = retime_s1_107_reg_reg_IQ;
 reg retime_s1_108_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_108_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_108_reg_reg_IQ <= mul_22_25_n_2108;
     end
 assign n_61 = retime_s1_108_reg_reg_IQ;
 reg retime_s1_109_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_109_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_109_reg_reg_IQ <= mul_22_25_n_2123;
     end
 assign n_60 = retime_s1_109_reg_reg_IQ;
 reg retime_s1_110_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_110_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_110_reg_reg_IQ <= mul_22_25_n_1684;
     end
 assign n_59 = retime_s1_110_reg_reg_IQ;
 reg retime_s1_111_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_111_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_111_reg_reg_IQ <= mul_22_25_n_1686;
     end
 assign n_58 = retime_s1_111_reg_reg_IQ;
 reg retime_s1_112_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_112_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_112_reg_reg_IQ <= mul_22_25_n_1255;
     end
 assign n_57 = retime_s1_112_reg_reg_IQ;
 reg retime_s1_113_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_113_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_113_reg_reg_IQ <= mul_22_25_n_1223;
     end
 assign n_56 = retime_s1_113_reg_reg_IQ;
 reg retime_s1_114_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_114_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_114_reg_reg_IQ <= mul_22_25_n_1253;
     end
 assign n_55 = retime_s1_114_reg_reg_IQ;
 reg retime_s1_115_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_115_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_115_reg_reg_IQ <= mul_22_25_n_1254;
     end
 assign n_54 = retime_s1_115_reg_reg_IQ;
 reg retime_s1_116_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_116_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_116_reg_reg_IQ <= mul_22_25_n_1608;
     end
 assign n_52 = retime_s1_116_reg_reg_IQ;
 reg retime_s1_117_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_117_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_117_reg_reg_IQ <= mul_22_25_n_1626;
     end
 assign n_51 = retime_s1_117_reg_reg_IQ;
 reg retime_s1_118_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_118_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_118_reg_reg_IQ <= mul_22_25_n_1539;
     end
 assign n_50 = retime_s1_118_reg_reg_IQ;
 reg retime_s1_119_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_119_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_119_reg_reg_IQ <= mul_22_25_n_1729;
     end
 assign n_49 = retime_s1_119_reg_reg_IQ;
 reg retime_s1_120_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_120_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_120_reg_reg_IQ <= mul_22_25_n_1752;
     end
 assign n_48 = retime_s1_120_reg_reg_IQ;
 reg retime_s1_121_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_121_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_121_reg_reg_IQ <= mul_22_25_n_1251;
     end
 assign n_47 = retime_s1_121_reg_reg_IQ;
 reg retime_s1_122_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_122_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_122_reg_reg_IQ <= mul_22_25_n_1538;
     end
 assign n_46 = retime_s1_122_reg_reg_IQ;
 reg retime_s1_123_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_123_reg_reg_IQ <= 1'B0;
     else begin
         retime_s1_123_reg_reg_IQ <= mul_22_25_n_1551;
     end
 assign n_45 = retime_s1_123_reg_reg_IQ;
 reg retime_s1_124_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_124_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_124_reg_reg_IQ <= mul_22_25_n_2090;
     end
 assign n_44 = retime_s1_124_reg_reg_IQ;
 reg retime_s1_125_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) retime_s1_125_reg_reg_IQ <= 1'B1;
     else begin
         retime_s1_125_reg_reg_IQ <= mul_22_25_n_2106;
     end
 assign n_43 = retime_s1_125_reg_reg_IQ;
 assign mul_22_25_n_1526 = ((mul_22_25_n_879 & mul_22_25_n_628) | (mul_22_25_n_644 & (mul_22_25_n_879
    ^ mul_22_25_n_628)));
 assign mul_22_25_n_1525 = (mul_22_25_n_644 ^ (mul_22_25_n_879 ^ mul_22_25_n_628));
 assign mul_22_25_n_2265 = ((mul_22_25_n_1066 & mul_22_25_n_906) | (mul_22_25_n_1162 & (mul_22_25_n_1066
    ^ mul_22_25_n_906)));
 assign mul_22_25_n_1524 = (mul_22_25_n_1162 ^ (mul_22_25_n_1066 ^ mul_22_25_n_906));
 assign mul_22_25_n_2224 = ((mul_22_25_n_655 & mul_22_25_n_624) | (mul_22_25_n_792 & (mul_22_25_n_655
    ^ mul_22_25_n_624)));
 assign mul_22_25_n_2225 = (mul_22_25_n_792 ^ (mul_22_25_n_655 ^ mul_22_25_n_624));
 assign mul_22_25_n_1523 = ((mul_22_25_n_1156 & mul_22_25_n_1017) | (mul_22_25_n_2225 & (mul_22_25_n_1156
    ^ mul_22_25_n_1017)));
 assign mul_22_25_n_1522 = (mul_22_25_n_2225 ^ (mul_22_25_n_1156 ^ mul_22_25_n_1017));
 assign mul_22_25_n_2222 = ((mul_22_25_n_779 & mul_22_25_n_1063) | (mul_22_25_n_773 & (mul_22_25_n_779
    ^ mul_22_25_n_1063)));
 assign mul_22_25_n_2223 = (mul_22_25_n_773 ^ (mul_22_25_n_779 ^ mul_22_25_n_1063));
 assign mul_22_25_n_1521 = ((mul_22_25_n_2224 & mul_22_25_n_1163) | (mul_22_25_n_2223 & (mul_22_25_n_2224
    ^ mul_22_25_n_1163)));
 assign mul_22_25_n_1520 = (mul_22_25_n_2223 ^ (mul_22_25_n_2224 ^ mul_22_25_n_1163));
 assign mul_22_25_n_2219 = ((mul_22_25_n_656 & mul_22_25_n_626) | (mul_22_25_n_829 & (mul_22_25_n_656
    ^ mul_22_25_n_626)));
 assign mul_22_25_n_2221 = (mul_22_25_n_829 ^ (mul_22_25_n_656 ^ mul_22_25_n_626));
 assign mul_22_25_n_2217 = ((mul_22_25_n_723 & mul_22_25_n_714) | (mul_22_25_n_1159 & (mul_22_25_n_723
    ^ mul_22_25_n_714)));
 assign mul_22_25_n_2220 = (mul_22_25_n_1159 ^ (mul_22_25_n_723 ^ mul_22_25_n_714));
 assign mul_22_25_n_2266 = ((mul_22_25_n_2221 & mul_22_25_n_2222) | (mul_22_25_n_2220 & (mul_22_25_n_2221
    ^ mul_22_25_n_2222)));
 assign mul_22_25_n_1519 = (mul_22_25_n_2220 ^ (mul_22_25_n_2221 ^ mul_22_25_n_2222));
 assign mul_22_25_n_2215 = ((mul_22_25_n_1062 & mul_22_25_n_705) | (mul_22_25_n_665 & (mul_22_25_n_1062
    ^ mul_22_25_n_705)));
 assign mul_22_25_n_2218 = (mul_22_25_n_665 ^ (mul_22_25_n_1062 ^ mul_22_25_n_705));
 assign mul_22_25_n_2212 = ((mul_22_25_n_1171 & mul_22_25_n_753) | (mul_22_25_n_2219 & (mul_22_25_n_1171
    ^ mul_22_25_n_753)));
 assign mul_22_25_n_2216 = (mul_22_25_n_2219 ^ (mul_22_25_n_1171 ^ mul_22_25_n_753));
 assign mul_22_25_n_1518 = ((mul_22_25_n_2217 & mul_22_25_n_2218) | (mul_22_25_n_2216 & (mul_22_25_n_2217
    ^ mul_22_25_n_2218)));
 assign mul_22_25_n_2226 = (mul_22_25_n_2216 ^ (mul_22_25_n_2217 ^ mul_22_25_n_2218));
 assign mul_22_25_n_2210 = ((mul_22_25_n_838 & mul_22_25_n_632) | (mul_22_25_n_747 & (mul_22_25_n_838
    ^ mul_22_25_n_632)));
 assign mul_22_25_n_2214 = (mul_22_25_n_747 ^ (mul_22_25_n_838 ^ mul_22_25_n_632));
 assign mul_22_25_n_2209 = ((mul_22_25_n_650 & mul_22_25_n_869) | (mul_22_25_n_988 & (mul_22_25_n_650
    ^ mul_22_25_n_869)));
 assign mul_22_25_n_2213 = (mul_22_25_n_988 ^ (mul_22_25_n_650 ^ mul_22_25_n_869));
 assign mul_22_25_n_2205 = ((mul_22_25_n_2215 & mul_22_25_n_1146) | (mul_22_25_n_2214 & (mul_22_25_n_2215
    ^ mul_22_25_n_1146)));
 assign mul_22_25_n_2211 = (mul_22_25_n_2214 ^ (mul_22_25_n_2215 ^ mul_22_25_n_1146));
 assign mul_22_25_n_1517 = ((mul_22_25_n_2212 & mul_22_25_n_2213) | (mul_22_25_n_2211 & (mul_22_25_n_2212
    ^ mul_22_25_n_2213)));
 assign mul_22_25_n_2227 = (mul_22_25_n_2211 ^ (mul_22_25_n_2212 ^ mul_22_25_n_2213));
 assign mul_22_25_n_2204 = ((mul_22_25_n_846 & mul_22_25_n_953) | (mul_22_25_n_649 & (mul_22_25_n_846
    ^ mul_22_25_n_953)));
 assign mul_22_25_n_2208 = (mul_22_25_n_649 ^ (mul_22_25_n_846 ^ mul_22_25_n_953));
 assign mul_22_25_n_2201 = ((mul_22_25_n_962 & mul_22_25_n_1068) | (mul_22_25_n_1174 & (mul_22_25_n_962
    ^ mul_22_25_n_1068)));
 assign mul_22_25_n_2207 = (mul_22_25_n_1174 ^ (mul_22_25_n_962 ^ mul_22_25_n_1068));
 assign mul_22_25_n_2199 = ((mul_22_25_n_2209 & mul_22_25_n_2210) | (mul_22_25_n_2208 & (mul_22_25_n_2209
    ^ mul_22_25_n_2210)));
 assign mul_22_25_n_2206 = (mul_22_25_n_2208 ^ (mul_22_25_n_2209 ^ mul_22_25_n_2210));
 assign mul_22_25_n_1516 = ((mul_22_25_n_2206 & mul_22_25_n_2207) | (mul_22_25_n_2205 & (mul_22_25_n_2206
    ^ mul_22_25_n_2207)));
 assign mul_22_25_n_1515 = (mul_22_25_n_2205 ^ (mul_22_25_n_2206 ^ mul_22_25_n_2207));
 assign mul_22_25_n_2197 = ((mul_22_25_n_939 & mul_22_25_n_634) | (mul_22_25_n_934 & (mul_22_25_n_939
    ^ mul_22_25_n_634)));
 assign mul_22_25_n_2202 = (mul_22_25_n_934 ^ (mul_22_25_n_939 ^ mul_22_25_n_634));
 assign mul_22_25_n_2196 = ((mul_22_25_n_648 & mul_22_25_n_923) | (mul_22_25_n_917 & (mul_22_25_n_648
    ^ mul_22_25_n_923)));
 assign mul_22_25_n_2203 = (mul_22_25_n_917 ^ (mul_22_25_n_648 ^ mul_22_25_n_923));
 assign mul_22_25_n_2193 = ((mul_22_25_n_1145 & mul_22_25_n_1092) | (mul_22_25_n_2204 & (mul_22_25_n_1145
    ^ mul_22_25_n_1092)));
 assign mul_22_25_n_2200 = (mul_22_25_n_2204 ^ (mul_22_25_n_1145 ^ mul_22_25_n_1092));
 assign mul_22_25_n_2191 = ((mul_22_25_n_2202 & mul_22_25_n_2203) | (mul_22_25_n_2201 & (mul_22_25_n_2202
    ^ mul_22_25_n_2203)));
 assign mul_22_25_n_2198 = (mul_22_25_n_2201 ^ (mul_22_25_n_2202 ^ mul_22_25_n_2203));
 assign mul_22_25_n_2267 = ((mul_22_25_n_2199 & mul_22_25_n_2200) | (mul_22_25_n_2198 & (mul_22_25_n_2199
    ^ mul_22_25_n_2200)));
 assign mul_22_25_n_1514 = (mul_22_25_n_2198 ^ (mul_22_25_n_2199 ^ mul_22_25_n_2200));
 assign mul_22_25_n_2189 = ((mul_22_25_n_902 & mul_22_25_n_812) | (mul_22_25_n_897 & (mul_22_25_n_902
    ^ mul_22_25_n_812)));
 assign mul_22_25_n_2194 = (mul_22_25_n_897 ^ (mul_22_25_n_902 ^ mul_22_25_n_812));
 assign mul_22_25_n_2188 = ((mul_22_25_n_886 & mul_22_25_n_890) | (mul_22_25_n_1060 & (mul_22_25_n_886
    ^ mul_22_25_n_890)));
 assign mul_22_25_n_2195 = (mul_22_25_n_1060 ^ (mul_22_25_n_886 ^ mul_22_25_n_890));
 assign mul_22_25_n_2184 = ((mul_22_25_n_2197 & mul_22_25_n_1166) | (mul_22_25_n_2196 & (mul_22_25_n_2197
    ^ mul_22_25_n_1166)));
 assign mul_22_25_n_2192 = (mul_22_25_n_2196 ^ (mul_22_25_n_2197 ^ mul_22_25_n_1166));
 assign mul_22_25_n_2181 = ((mul_22_25_n_2194 & mul_22_25_n_2195) | (mul_22_25_n_2193 & (mul_22_25_n_2194
    ^ mul_22_25_n_2195)));
 assign mul_22_25_n_2190 = (mul_22_25_n_2193 ^ (mul_22_25_n_2194 ^ mul_22_25_n_2195));
 assign mul_22_25_n_2268 = ((mul_22_25_n_2191 & mul_22_25_n_2192) | (mul_22_25_n_2190 & (mul_22_25_n_2191
    ^ mul_22_25_n_2192)));
 assign mul_22_25_n_2228 = (mul_22_25_n_2190 ^ (mul_22_25_n_2191 ^ mul_22_25_n_2192));
 assign mul_22_25_n_2180 = ((mul_22_25_n_643 & mul_22_25_n_627) | (mul_22_25_n_841 & (mul_22_25_n_643
    ^ mul_22_25_n_627)));
 assign mul_22_25_n_2187 = (mul_22_25_n_841 ^ (mul_22_25_n_643 ^ mul_22_25_n_627));
 assign mul_22_25_n_2179 = ((mul_22_25_n_827 & mul_22_25_n_832) | (mul_22_25_n_981 & (mul_22_25_n_827
    ^ mul_22_25_n_832)));
 assign mul_22_25_n_2186 = (mul_22_25_n_981 ^ (mul_22_25_n_827 ^ mul_22_25_n_832));
 assign mul_22_25_n_2176 = ((mul_22_25_n_750 & mul_22_25_n_813) | (mul_22_25_n_1157 & (mul_22_25_n_750
    ^ mul_22_25_n_813)));
 assign mul_22_25_n_2185 = (mul_22_25_n_1157 ^ (mul_22_25_n_750 ^ mul_22_25_n_813));
 assign mul_22_25_n_2174 = ((mul_22_25_n_2188 & mul_22_25_n_2189) | (mul_22_25_n_2187 & (mul_22_25_n_2188
    ^ mul_22_25_n_2189)));
 assign mul_22_25_n_2183 = (mul_22_25_n_2187 ^ (mul_22_25_n_2188 ^ mul_22_25_n_2189));
 assign mul_22_25_n_2172 = ((mul_22_25_n_2185 & mul_22_25_n_2186) | (mul_22_25_n_2184 & (mul_22_25_n_2185
    ^ mul_22_25_n_2186)));
 assign mul_22_25_n_2182 = (mul_22_25_n_2184 ^ (mul_22_25_n_2185 ^ mul_22_25_n_2186));
 assign mul_22_25_n_2269 = ((mul_22_25_n_2182 & mul_22_25_n_2183) | (mul_22_25_n_2181 & (mul_22_25_n_2182
    ^ mul_22_25_n_2183)));
 assign mul_22_25_n_2229 = (mul_22_25_n_2181 ^ (mul_22_25_n_2182 ^ mul_22_25_n_2183));
 assign mul_22_25_n_2170 = ((mul_22_25_n_1064 & mul_22_25_n_845) | (mul_22_25_n_791 & (mul_22_25_n_1064
    ^ mul_22_25_n_845)));
 assign mul_22_25_n_2177 = (mul_22_25_n_791 ^ (mul_22_25_n_1064 ^ mul_22_25_n_845));
 assign mul_22_25_n_2169 = ((mul_22_25_n_950 & mul_22_25_n_786) | (mul_22_25_n_870 & (mul_22_25_n_950
    ^ mul_22_25_n_786)));
 assign mul_22_25_n_2178 = (mul_22_25_n_870 ^ (mul_22_25_n_950 ^ mul_22_25_n_786));
 assign mul_22_25_n_2165 = ((mul_22_25_n_1168 & mul_22_25_n_771) | (mul_22_25_n_2180 & (mul_22_25_n_1168
    ^ mul_22_25_n_771)));
 assign mul_22_25_n_2175 = (mul_22_25_n_2180 ^ (mul_22_25_n_1168 ^ mul_22_25_n_771));
 assign mul_22_25_n_2163 = ((mul_22_25_n_2178 & mul_22_25_n_2179) | (mul_22_25_n_2177 & (mul_22_25_n_2178
    ^ mul_22_25_n_2179)));
 assign mul_22_25_n_2173 = (mul_22_25_n_2177 ^ (mul_22_25_n_2178 ^ mul_22_25_n_2179));
 assign mul_22_25_n_2161 = ((mul_22_25_n_2175 & mul_22_25_n_2176) | (mul_22_25_n_2174 & (mul_22_25_n_2175
    ^ mul_22_25_n_2176)));
 assign mul_22_25_n_2171 = (mul_22_25_n_2174 ^ (mul_22_25_n_2175 ^ mul_22_25_n_2176));
 assign mul_22_25_n_2270 = ((mul_22_25_n_2172 & mul_22_25_n_2173) | (mul_22_25_n_2171 & (mul_22_25_n_2172
    ^ mul_22_25_n_2173)));
 assign mul_22_25_n_2230 = (mul_22_25_n_2171 ^ (mul_22_25_n_2172 ^ mul_22_25_n_2173));
 assign mul_22_25_n_2159 = ((mul_22_25_n_642 & mul_22_25_n_630) | (mul_22_25_n_749 & (mul_22_25_n_642
    ^ mul_22_25_n_630)));
 assign mul_22_25_n_2167 = (mul_22_25_n_749 ^ (mul_22_25_n_642 ^ mul_22_25_n_630));
 assign mul_22_25_n_2157 = ((mul_22_25_n_738 & mul_22_25_n_740) | (mul_22_25_n_722 & (mul_22_25_n_738
    ^ mul_22_25_n_740)));
 assign mul_22_25_n_2166 = (mul_22_25_n_722 ^ (mul_22_25_n_738 ^ mul_22_25_n_740));
 assign mul_22_25_n_2158 = ((mul_22_25_n_697 & mul_22_25_n_1019) | (mul_22_25_n_726 & (mul_22_25_n_697
    ^ mul_22_25_n_1019)));
 assign mul_22_25_n_2168 = (mul_22_25_n_726 ^ (mul_22_25_n_697 ^ mul_22_25_n_1019));
 assign mul_22_25_n_2153 = ((mul_22_25_n_2170 & mul_22_25_n_1155) | (mul_22_25_n_2169 & (mul_22_25_n_2170
    ^ mul_22_25_n_1155)));
 assign mul_22_25_n_2164 = (mul_22_25_n_2169 ^ (mul_22_25_n_2170 ^ mul_22_25_n_1155));
 assign mul_22_25_n_2151 = ((mul_22_25_n_2167 & mul_22_25_n_2168) | (mul_22_25_n_2166 & (mul_22_25_n_2167
    ^ mul_22_25_n_2168)));
 assign mul_22_25_n_2162 = (mul_22_25_n_2166 ^ (mul_22_25_n_2167 ^ mul_22_25_n_2168));
 assign mul_22_25_n_2149 = ((mul_22_25_n_2164 & mul_22_25_n_2165) | (mul_22_25_n_2163 & (mul_22_25_n_2164
    ^ mul_22_25_n_2165)));
 assign mul_22_25_n_2160 = (mul_22_25_n_2163 ^ (mul_22_25_n_2164 ^ mul_22_25_n_2165));
 assign mul_22_25_n_2271 = ((mul_22_25_n_2161 & mul_22_25_n_2162) | (mul_22_25_n_2160 & (mul_22_25_n_2161
    ^ mul_22_25_n_2162)));
 assign mul_22_25_n_2231 = (mul_22_25_n_2160 ^ (mul_22_25_n_2161 ^ mul_22_25_n_2162));
 assign mul_22_25_n_2147 = ((mul_22_25_n_702 & mul_22_25_n_704) | (mul_22_25_n_1061 & (mul_22_25_n_702
    ^ mul_22_25_n_704)));
 assign mul_22_25_n_2156 = (mul_22_25_n_1061 ^ (mul_22_25_n_702 ^ mul_22_25_n_704));
 assign mul_22_25_n_2146 = ((mul_22_25_n_695 & mul_22_25_n_918) | (mul_22_25_n_970 & (mul_22_25_n_695
    ^ mul_22_25_n_918)));
 assign mul_22_25_n_2155 = (mul_22_25_n_970 ^ (mul_22_25_n_695 ^ mul_22_25_n_918));
 assign mul_22_25_n_2142 = ((mul_22_25_n_1009 & mul_22_25_n_866) | (mul_22_25_n_1164 & (mul_22_25_n_1009
    ^ mul_22_25_n_866)));
 assign mul_22_25_n_2154 = (mul_22_25_n_1164 ^ (mul_22_25_n_1009 ^ mul_22_25_n_866));
 assign mul_22_25_n_2140 = ((mul_22_25_n_2158 & mul_22_25_n_2159) | (mul_22_25_n_2157 & (mul_22_25_n_2158
    ^ mul_22_25_n_2159)));
 assign mul_22_25_n_2152 = (mul_22_25_n_2157 ^ (mul_22_25_n_2158 ^ mul_22_25_n_2159));
 assign mul_22_25_n_2139 = ((mul_22_25_n_2155 & mul_22_25_n_2156) | (mul_22_25_n_2154 & (mul_22_25_n_2155
    ^ mul_22_25_n_2156)));
 assign mul_22_25_n_2150 = (mul_22_25_n_2154 ^ (mul_22_25_n_2155 ^ mul_22_25_n_2156));
 assign mul_22_25_n_2136 = ((mul_22_25_n_2152 & mul_22_25_n_2153) | (mul_22_25_n_2151 & (mul_22_25_n_2152
    ^ mul_22_25_n_2153)));
 assign mul_22_25_n_2148 = (mul_22_25_n_2151 ^ (mul_22_25_n_2152 ^ mul_22_25_n_2153));
 assign mul_22_25_n_2272 = ((mul_22_25_n_2149 & mul_22_25_n_2150) | (mul_22_25_n_2148 & (mul_22_25_n_2149
    ^ mul_22_25_n_2150)));
 assign mul_22_25_n_2232 = (mul_22_25_n_2148 ^ (mul_22_25_n_2149 ^ mul_22_25_n_2150));
 assign mul_22_25_n_2134 = ((mul_22_25_n_666 & mul_22_25_n_635) | (mul_22_25_n_833 & (mul_22_25_n_666
    ^ mul_22_25_n_635)));
 assign mul_22_25_n_2144 = (mul_22_25_n_833 ^ (mul_22_25_n_666 ^ mul_22_25_n_635));
 assign mul_22_25_n_2133 = ((mul_22_25_n_835 & mul_22_25_n_801) | (mul_22_25_n_1020 & (mul_22_25_n_835
    ^ mul_22_25_n_801)));
 assign mul_22_25_n_2143 = (mul_22_25_n_1020 ^ (mul_22_25_n_835 ^ mul_22_25_n_801));
 assign mul_22_25_n_2132 = ((mul_22_25_n_1011 & mul_22_25_n_907) | (mul_22_25_n_784 & (mul_22_25_n_1011
    ^ mul_22_25_n_907)));
 assign mul_22_25_n_2145 = (mul_22_25_n_784 ^ (mul_22_25_n_1011 ^ mul_22_25_n_907));
 assign mul_22_25_n_2128 = ((mul_22_25_n_1154 & mul_22_25_n_861) | (mul_22_25_n_2147 & (mul_22_25_n_1154
    ^ mul_22_25_n_861)));
 assign mul_22_25_n_2141 = (mul_22_25_n_2147 ^ (mul_22_25_n_1154 ^ mul_22_25_n_861));
 assign mul_22_25_n_2126 = ((mul_22_25_n_2145 & mul_22_25_n_2146) | (mul_22_25_n_2144 & (mul_22_25_n_2145
    ^ mul_22_25_n_2146)));
 assign mul_22_25_n_2138 = (mul_22_25_n_2144 ^ (mul_22_25_n_2145 ^ mul_22_25_n_2146));
 assign mul_22_25_n_2124 = ((mul_22_25_n_2142 & mul_22_25_n_2143) | (mul_22_25_n_2141 & (mul_22_25_n_2142
    ^ mul_22_25_n_2143)));
 assign mul_22_25_n_2137 = (mul_22_25_n_2141 ^ (mul_22_25_n_2142 ^ mul_22_25_n_2143));
 assign mul_22_25_n_2122 = ((mul_22_25_n_2139 & mul_22_25_n_2140) | (mul_22_25_n_2138 & (mul_22_25_n_2139
    ^ mul_22_25_n_2140)));
 assign mul_22_25_n_2135 = (mul_22_25_n_2138 ^ (mul_22_25_n_2139 ^ mul_22_25_n_2140));
 assign mul_22_25_n_2273 = ((mul_22_25_n_2136 & mul_22_25_n_2137) | (mul_22_25_n_2135 & (mul_22_25_n_2136
    ^ mul_22_25_n_2137)));
 assign mul_22_25_n_2233 = (mul_22_25_n_2135 ^ (mul_22_25_n_2136 ^ mul_22_25_n_2137));
 assign mul_22_25_n_2120 = ((mul_22_25_n_928 & mul_22_25_n_987) | (mul_22_25_n_888 & (mul_22_25_n_928
    ^ mul_22_25_n_987)));
 assign mul_22_25_n_2130 = (mul_22_25_n_888 ^ (mul_22_25_n_928 ^ mul_22_25_n_987));
 assign mul_22_25_n_2118 = ((mul_22_25_n_1067 & mul_22_25_n_896) | (mul_22_25_n_1015 & (mul_22_25_n_1067
    ^ mul_22_25_n_896)));
 assign mul_22_25_n_2129 = (mul_22_25_n_1015 ^ (mul_22_25_n_1067 ^ mul_22_25_n_896));
 assign mul_22_25_n_2119 = ((mul_22_25_n_967 & mul_22_25_n_969) | (mul_22_25_n_905 & (mul_22_25_n_967
    ^ mul_22_25_n_969)));
 assign mul_22_25_n_2131 = (mul_22_25_n_905 ^ (mul_22_25_n_967 ^ mul_22_25_n_969));
 assign mul_22_25_n_2113 = ((mul_22_25_n_2134 & mul_22_25_n_1167) | (mul_22_25_n_2133 & (mul_22_25_n_2134
    ^ mul_22_25_n_1167)));
 assign mul_22_25_n_2127 = (mul_22_25_n_2133 ^ (mul_22_25_n_2134 ^ mul_22_25_n_1167));
 assign mul_22_25_n_2112 = ((mul_22_25_n_2131 & mul_22_25_n_2132) | (mul_22_25_n_2130 & (mul_22_25_n_2131
    ^ mul_22_25_n_2132)));
 assign mul_22_25_n_2125 = (mul_22_25_n_2130 ^ (mul_22_25_n_2131 ^ mul_22_25_n_2132));
 assign mul_22_25_n_2108 = ((mul_22_25_n_2128 & mul_22_25_n_2129) | (mul_22_25_n_2127 & (mul_22_25_n_2128
    ^ mul_22_25_n_2129)));
 assign mul_22_25_n_2123 = (mul_22_25_n_2127 ^ (mul_22_25_n_2128 ^ mul_22_25_n_2129));
 assign mul_22_25_n_2107 = ((mul_22_25_n_2125 & mul_22_25_n_2126) | (mul_22_25_n_2124 & (mul_22_25_n_2125
    ^ mul_22_25_n_2126)));
 assign mul_22_25_n_2121 = (mul_22_25_n_2124 ^ (mul_22_25_n_2125 ^ mul_22_25_n_2126));
 assign mul_22_25_n_2274 = ((n_92 & n_60) | (n_66 & (n_92 ^ n_60)));
 assign mul_22_25_n_2234 = (n_66 ^ (n_92 ^ n_60));
 assign mul_22_25_n_2104 = ((mul_22_25_n_647 & mul_22_25_n_629) | (mul_22_25_n_946 & (mul_22_25_n_647
    ^ mul_22_25_n_629)));
 assign mul_22_25_n_2117 = (mul_22_25_n_946 ^ (mul_22_25_n_647 ^ mul_22_25_n_629));
 assign mul_22_25_n_2105 = ((mul_22_25_n_1050 & mul_22_25_n_942) | (mul_22_25_n_938 & (mul_22_25_n_1050
    ^ mul_22_25_n_942)));
 assign mul_22_25_n_2116 = (mul_22_25_n_938 ^ (mul_22_25_n_1050 ^ mul_22_25_n_942));
 assign mul_22_25_n_2103 = ((mul_22_25_n_930 & mul_22_25_n_932) | (mul_22_25_n_729 & (mul_22_25_n_930
    ^ mul_22_25_n_932)));
 assign mul_22_25_n_2115 = (mul_22_25_n_729 ^ (mul_22_25_n_930 ^ mul_22_25_n_932));
 assign mul_22_25_n_2099 = ((mul_22_25_n_922 & mul_22_25_n_924) | (mul_22_25_n_1158 & (mul_22_25_n_922
    ^ mul_22_25_n_924)));
 assign mul_22_25_n_2114 = (mul_22_25_n_1158 ^ (mul_22_25_n_922 ^ mul_22_25_n_924));
 assign mul_22_25_n_2098 = ((mul_22_25_n_2119 & mul_22_25_n_2120) | (mul_22_25_n_2118 & (mul_22_25_n_2119
    ^ mul_22_25_n_2120)));
 assign mul_22_25_n_2111 = (mul_22_25_n_2118 ^ (mul_22_25_n_2119 ^ mul_22_25_n_2120));
 assign mul_22_25_n_2095 = ((mul_22_25_n_2116 & mul_22_25_n_2117) | (mul_22_25_n_2115 & (mul_22_25_n_2116
    ^ mul_22_25_n_2117)));
 assign mul_22_25_n_2110 = (mul_22_25_n_2115 ^ (mul_22_25_n_2116 ^ mul_22_25_n_2117));
 assign mul_22_25_n_2092 = ((mul_22_25_n_2113 & mul_22_25_n_2114) | (mul_22_25_n_2112 & (mul_22_25_n_2113
    ^ mul_22_25_n_2114)));
 assign mul_22_25_n_2109 = (mul_22_25_n_2112 ^ (mul_22_25_n_2113 ^ mul_22_25_n_2114));
 assign mul_22_25_n_2090 = ((mul_22_25_n_2110 & mul_22_25_n_2111) | (mul_22_25_n_2109 & (mul_22_25_n_2110
    ^ mul_22_25_n_2111)));
 assign mul_22_25_n_2106 = (mul_22_25_n_2109 ^ (mul_22_25_n_2110 ^ mul_22_25_n_2111));
 assign mul_22_25_n_2275 = ((n_67 & n_61) | (n_43 & (n_67 ^ n_61)));
 assign mul_22_25_n_2235 = (n_43 ^ (n_67 ^ n_61));
 assign mul_22_25_n_2087 = ((mul_22_25_n_1105 & mul_22_25_n_1103) | (mul_22_25_n_1109 & (mul_22_25_n_1105
    ^ mul_22_25_n_1103)));
 assign mul_22_25_n_2101 = (mul_22_25_n_1109 ^ (mul_22_25_n_1105 ^ mul_22_25_n_1103));
 assign mul_22_25_n_2088 = ((mul_22_25_n_768 & mul_22_25_n_721) | (mul_22_25_n_1058 & (mul_22_25_n_768
    ^ mul_22_25_n_721)));
 assign mul_22_25_n_2100 = (mul_22_25_n_1058 ^ (mul_22_25_n_768 ^ mul_22_25_n_721));
 assign mul_22_25_n_2089 = ((mul_22_25_n_903 & mul_22_25_n_645) | (mul_22_25_n_899 & (mul_22_25_n_903
    ^ mul_22_25_n_645)));
 assign mul_22_25_n_2102 = (mul_22_25_n_899 ^ (mul_22_25_n_903 ^ mul_22_25_n_645));
 assign mul_22_25_n_2082 = ((mul_22_25_n_1172 & mul_22_25_n_920) | (mul_22_25_n_2105 & (mul_22_25_n_1172
    ^ mul_22_25_n_920)));
 assign mul_22_25_n_2097 = (mul_22_25_n_2105 ^ (mul_22_25_n_1172 ^ mul_22_25_n_920));
 assign mul_22_25_n_2081 = ((mul_22_25_n_2103 & mul_22_25_n_2104) | (mul_22_25_n_2102 & (mul_22_25_n_2103
    ^ mul_22_25_n_2104)));
 assign mul_22_25_n_2096 = (mul_22_25_n_2102 ^ (mul_22_25_n_2103 ^ mul_22_25_n_2104));
 assign mul_22_25_n_2079 = ((mul_22_25_n_2100 & mul_22_25_n_2101) | (mul_22_25_n_2099 & (mul_22_25_n_2100
    ^ mul_22_25_n_2101)));
 assign mul_22_25_n_2094 = (mul_22_25_n_2099 ^ (mul_22_25_n_2100 ^ mul_22_25_n_2101));
 assign mul_22_25_n_2076 = ((mul_22_25_n_2097 & mul_22_25_n_2098) | (mul_22_25_n_2096 & (mul_22_25_n_2097
    ^ mul_22_25_n_2098)));
 assign mul_22_25_n_2093 = (mul_22_25_n_2096 ^ (mul_22_25_n_2097 ^ mul_22_25_n_2098));
 assign mul_22_25_n_2073 = ((mul_22_25_n_2094 & mul_22_25_n_2095) | (mul_22_25_n_2093 & (mul_22_25_n_2094
    ^ mul_22_25_n_2095)));
 assign mul_22_25_n_2091 = (mul_22_25_n_2093 ^ (mul_22_25_n_2094 ^ mul_22_25_n_2095));
 assign mul_22_25_n_2276 = ((n_152 & n_161) | (n_44 & (n_152 ^ n_161)));
 assign mul_22_25_n_2236 = (n_44 ^ (n_152 ^ n_161));
 assign mul_22_25_n_2070 = ((mul_22_25_n_867 & mul_22_25_n_625) | (mul_22_25_n_864 & (mul_22_25_n_867
    ^ mul_22_25_n_625)));
 assign mul_22_25_n_2083 = (mul_22_25_n_864 ^ (mul_22_25_n_867 ^ mul_22_25_n_625));
 assign mul_22_25_n_2069 = ((mul_22_25_n_871 & mul_22_25_n_859) | (mul_22_25_n_858 & (mul_22_25_n_871
    ^ mul_22_25_n_859)));
 assign mul_22_25_n_2085 = (mul_22_25_n_858 ^ (mul_22_25_n_871 ^ mul_22_25_n_859));
 assign mul_22_25_n_2072 = ((mul_22_25_n_959 & mul_22_25_n_854) | (mul_22_25_n_653 & (mul_22_25_n_959
    ^ mul_22_25_n_854)));
 assign mul_22_25_n_2084 = (mul_22_25_n_653 ^ (mul_22_25_n_959 ^ mul_22_25_n_854));
 assign mul_22_25_n_2071 = ((mul_22_25_n_844 & mul_22_25_n_849) | (mul_22_25_n_843 & (mul_22_25_n_844
    ^ mul_22_25_n_849)));
 assign mul_22_25_n_2086 = (mul_22_25_n_843 ^ (mul_22_25_n_844 ^ mul_22_25_n_849));
 assign mul_22_25_n_2064 = ((mul_22_25_n_2089 & mul_22_25_n_1147) | (mul_22_25_n_2088 & (mul_22_25_n_2089
    ^ mul_22_25_n_1147)));
 assign mul_22_25_n_2080 = (mul_22_25_n_2088 ^ (mul_22_25_n_2089 ^ mul_22_25_n_1147));
 assign mul_22_25_n_2062 = ((mul_22_25_n_2086 & mul_22_25_n_2087) | (mul_22_25_n_2085 & (mul_22_25_n_2086
    ^ mul_22_25_n_2087)));
 assign mul_22_25_n_2078 = (mul_22_25_n_2085 ^ (mul_22_25_n_2086 ^ mul_22_25_n_2087));
 assign mul_22_25_n_2059 = ((mul_22_25_n_2083 & mul_22_25_n_2084) | (mul_22_25_n_2082 & (mul_22_25_n_2083
    ^ mul_22_25_n_2084)));
 assign mul_22_25_n_2077 = (mul_22_25_n_2082 ^ (mul_22_25_n_2083 ^ mul_22_25_n_2084));
 assign mul_22_25_n_2057 = ((mul_22_25_n_2080 & mul_22_25_n_2081) | (mul_22_25_n_2079 & (mul_22_25_n_2080
    ^ mul_22_25_n_2081)));
 assign mul_22_25_n_2075 = (mul_22_25_n_2079 ^ (mul_22_25_n_2080 ^ mul_22_25_n_2081));
 assign mul_22_25_n_2056 = ((mul_22_25_n_2077 & mul_22_25_n_2078) | (mul_22_25_n_2076 & (mul_22_25_n_2077
    ^ mul_22_25_n_2078)));
 assign mul_22_25_n_2074 = (mul_22_25_n_2076 ^ (mul_22_25_n_2077 ^ mul_22_25_n_2078));
 assign mul_22_25_n_2277 = ((n_170 & n_150) | (n_153 & (n_170 ^ n_150)));
 assign mul_22_25_n_2237 = (n_153 ^ (n_170 ^ n_150));
 assign mul_22_25_n_2052 = ((mul_22_25_n_818 & mul_22_25_n_1055) | (mul_22_25_n_816 & (mul_22_25_n_818
    ^ mul_22_25_n_1055)));
 assign mul_22_25_n_2066 = (mul_22_25_n_816 ^ (mul_22_25_n_818 ^ mul_22_25_n_1055));
 assign mul_22_25_n_2054 = ((mul_22_25_n_810 & mul_22_25_n_752) | (mul_22_25_n_806 & (mul_22_25_n_810
    ^ mul_22_25_n_752)));
 assign mul_22_25_n_2067 = (mul_22_25_n_806 ^ (mul_22_25_n_810 ^ mul_22_25_n_752));
 assign mul_22_25_n_2053 = ((mul_22_25_n_837 & mul_22_25_n_641) | (mul_22_25_n_1057 & (mul_22_25_n_837
    ^ mul_22_25_n_641)));
 assign mul_22_25_n_2068 = (mul_22_25_n_1057 ^ (mul_22_25_n_837 ^ mul_22_25_n_641));
 assign mul_22_25_n_2047 = ((mul_22_25_n_803 & mul_22_25_n_694) | (mul_22_25_n_1175 & (mul_22_25_n_803
    ^ mul_22_25_n_694)));
 assign mul_22_25_n_2065 = (mul_22_25_n_1175 ^ (mul_22_25_n_803 ^ mul_22_25_n_694));
 assign mul_22_25_n_2046 = ((mul_22_25_n_2071 & mul_22_25_n_2072) | (mul_22_25_n_2070 & (mul_22_25_n_2071
    ^ mul_22_25_n_2072)));
 assign mul_22_25_n_2063 = (mul_22_25_n_2070 ^ (mul_22_25_n_2071 ^ mul_22_25_n_2072));
 assign mul_22_25_n_2043 = ((mul_22_25_n_2068 & mul_22_25_n_2069) | (mul_22_25_n_2067 & (mul_22_25_n_2068
    ^ mul_22_25_n_2069)));
 assign mul_22_25_n_2061 = (mul_22_25_n_2067 ^ (mul_22_25_n_2068 ^ mul_22_25_n_2069));
 assign mul_22_25_n_2041 = ((mul_22_25_n_2065 & mul_22_25_n_2066) | (mul_22_25_n_2064 & (mul_22_25_n_2065
    ^ mul_22_25_n_2066)));
 assign mul_22_25_n_2060 = (mul_22_25_n_2064 ^ (mul_22_25_n_2065 ^ mul_22_25_n_2066));
 assign mul_22_25_n_2039 = ((mul_22_25_n_2062 & mul_22_25_n_2063) | (mul_22_25_n_2061 & (mul_22_25_n_2062
    ^ mul_22_25_n_2063)));
 assign mul_22_25_n_2058 = (mul_22_25_n_2061 ^ (mul_22_25_n_2062 ^ mul_22_25_n_2063));
 assign mul_22_25_n_2036 = ((mul_22_25_n_2059 & mul_22_25_n_2060) | (mul_22_25_n_2058 & (mul_22_25_n_2059
    ^ mul_22_25_n_2060)));
 assign mul_22_25_n_2055 = (mul_22_25_n_2058 ^ (mul_22_25_n_2059 ^ mul_22_25_n_2060));
 assign mul_22_25_n_2278 = ((n_171 & n_151) | (n_144 & (n_171 ^ n_151)));
 assign mul_22_25_n_2238 = (n_144 ^ (n_171 ^ n_151));
 assign mul_22_25_n_2032 = ((mul_22_25_n_787 & mul_22_25_n_623) | (mul_22_25_n_785 & (mul_22_25_n_787
    ^ mul_22_25_n_623)));
 assign mul_22_25_n_2049 = (mul_22_25_n_785 ^ (mul_22_25_n_787 ^ mul_22_25_n_623));
 assign mul_22_25_n_2035 = ((mul_22_25_n_875 & mul_22_25_n_780) | (mul_22_25_n_776 & (mul_22_25_n_875
    ^ mul_22_25_n_780)));
 assign mul_22_25_n_2048 = (mul_22_25_n_776 ^ (mul_22_25_n_875 ^ mul_22_25_n_780));
 assign mul_22_25_n_2034 = ((mul_22_25_n_755 & mul_22_25_n_774) | (mul_22_25_n_683 & (mul_22_25_n_755
    ^ mul_22_25_n_774)));
 assign mul_22_25_n_2050 = (mul_22_25_n_683 ^ (mul_22_25_n_755 ^ mul_22_25_n_774));
 assign mul_22_25_n_2033 = ((mul_22_25_n_725 & mul_22_25_n_713) | (mul_22_25_n_758 & (mul_22_25_n_725
    ^ mul_22_25_n_713)));
 assign mul_22_25_n_2051 = (mul_22_25_n_758 ^ (mul_22_25_n_725 ^ mul_22_25_n_713));
 assign mul_22_25_n_2027 = ((mul_22_25_n_1148 & mul_22_25_n_766) | (mul_22_25_n_2054 & (mul_22_25_n_1148
    ^ mul_22_25_n_766)));
 assign mul_22_25_n_2045 = (mul_22_25_n_2054 ^ (mul_22_25_n_1148 ^ mul_22_25_n_766));
 assign mul_22_25_n_2024 = ((mul_22_25_n_2052 & mul_22_25_n_2053) | (mul_22_25_n_2051 & (mul_22_25_n_2052
    ^ mul_22_25_n_2053)));
 assign mul_22_25_n_2044 = (mul_22_25_n_2051 ^ (mul_22_25_n_2052 ^ mul_22_25_n_2053));
 assign mul_22_25_n_2025 = ((mul_22_25_n_2049 & mul_22_25_n_2050) | (mul_22_25_n_2048 & (mul_22_25_n_2049
    ^ mul_22_25_n_2050)));
 assign mul_22_25_n_2042 = (mul_22_25_n_2048 ^ (mul_22_25_n_2049 ^ mul_22_25_n_2050));
 assign mul_22_25_n_2021 = ((mul_22_25_n_2046 & mul_22_25_n_2047) | (mul_22_25_n_2045 & (mul_22_25_n_2046
    ^ mul_22_25_n_2047)));
 assign mul_22_25_n_2040 = (mul_22_25_n_2045 ^ (mul_22_25_n_2046 ^ mul_22_25_n_2047));
 assign mul_22_25_n_2020 = ((mul_22_25_n_2043 & mul_22_25_n_2044) | (mul_22_25_n_2042 & (mul_22_25_n_2043
    ^ mul_22_25_n_2044)));
 assign mul_22_25_n_2038 = (mul_22_25_n_2042 ^ (mul_22_25_n_2043 ^ mul_22_25_n_2044));
 assign mul_22_25_n_2017 = ((mul_22_25_n_2040 & mul_22_25_n_2041) | (mul_22_25_n_2039 & (mul_22_25_n_2040
    ^ mul_22_25_n_2041)));
 assign mul_22_25_n_2037 = (mul_22_25_n_2039 ^ (mul_22_25_n_2040 ^ mul_22_25_n_2041));
 assign mul_22_25_n_2279 = ((n_138 & n_157) | (n_145 & (n_138 ^ n_157)));
 assign mul_22_25_n_2239 = (n_145 ^ (n_138 ^ n_157));
 assign mul_22_25_n_2015 = ((mul_22_25_n_865 & mul_22_25_n_799) | (mul_22_25_n_748 & (mul_22_25_n_865
    ^ mul_22_25_n_799)));
 assign mul_22_25_n_2030 = (mul_22_25_n_748 ^ (mul_22_25_n_865 ^ mul_22_25_n_799));
 assign mul_22_25_n_2014 = ((mul_22_25_n_997 & mul_22_25_n_982) | (mul_22_25_n_925 & (mul_22_25_n_997
    ^ mul_22_25_n_982)));
 assign mul_22_25_n_2029 = (mul_22_25_n_925 ^ (mul_22_25_n_997 ^ mul_22_25_n_982));
 assign mul_22_25_n_2013 = ((mul_22_25_n_735 & mul_22_25_n_654) | (mul_22_25_n_733 & (mul_22_25_n_735
    ^ mul_22_25_n_654)));
 assign mul_22_25_n_2028 = (mul_22_25_n_733 ^ (mul_22_25_n_735 ^ mul_22_25_n_654));
 assign mul_22_25_n_2012 = ((mul_22_25_n_991 & mul_22_25_n_1059) | (mul_22_25_n_1027 & (mul_22_25_n_991
    ^ mul_22_25_n_1059)));
 assign mul_22_25_n_2031 = (mul_22_25_n_1027 ^ (mul_22_25_n_991 ^ mul_22_25_n_1059));
 assign mul_22_25_n_2006 = ((mul_22_25_n_2035 & mul_22_25_n_1170) | (mul_22_25_n_2034 & (mul_22_25_n_2035
    ^ mul_22_25_n_1170)));
 assign mul_22_25_n_2023 = (mul_22_25_n_2034 ^ (mul_22_25_n_2035 ^ mul_22_25_n_1170));
 assign mul_22_25_n_2005 = ((mul_22_25_n_2032 & mul_22_25_n_2033) | (mul_22_25_n_2031 & (mul_22_25_n_2032
    ^ mul_22_25_n_2033)));
 assign mul_22_25_n_2026 = (mul_22_25_n_2031 ^ (mul_22_25_n_2032 ^ mul_22_25_n_2033));
 assign mul_22_25_n_2004 = ((mul_22_25_n_2029 & mul_22_25_n_2030) | (mul_22_25_n_2028 & (mul_22_25_n_2029
    ^ mul_22_25_n_2030)));
 assign mul_22_25_n_2022 = (mul_22_25_n_2028 ^ (mul_22_25_n_2029 ^ mul_22_25_n_2030));
 assign mul_22_25_n_2000 = ((mul_22_25_n_2026 & mul_22_25_n_2027) | (mul_22_25_n_2025 & (mul_22_25_n_2026
    ^ mul_22_25_n_2027)));
 assign mul_22_25_n_2019 = (mul_22_25_n_2025 ^ (mul_22_25_n_2026 ^ mul_22_25_n_2027));
 assign mul_22_25_n_1998 = ((mul_22_25_n_2023 & mul_22_25_n_2024) | (mul_22_25_n_2022 & (mul_22_25_n_2023
    ^ mul_22_25_n_2024)));
 assign mul_22_25_n_2018 = (mul_22_25_n_2022 ^ (mul_22_25_n_2023 ^ mul_22_25_n_2024));
 assign mul_22_25_n_1996 = ((mul_22_25_n_2020 & mul_22_25_n_2021) | (mul_22_25_n_2019 & (mul_22_25_n_2020
    ^ mul_22_25_n_2021)));
 assign mul_22_25_n_2016 = (mul_22_25_n_2019 ^ (mul_22_25_n_2020 ^ mul_22_25_n_2021));
 assign mul_22_25_n_2280 = ((n_139 & n_166) | (n_71 & (n_139 ^ n_166)));
 assign mul_22_25_n_2240 = (n_71 ^ (n_139 ^ n_166));
 assign mul_22_25_n_1994 = ((mul_22_25_n_1005 & mul_22_25_n_631) | (mul_22_25_n_815 & (mul_22_25_n_1005
    ^ mul_22_25_n_631)));
 assign mul_22_25_n_2011 = (mul_22_25_n_815 ^ (mul_22_25_n_1005 ^ mul_22_25_n_631));
 assign mul_22_25_n_1993 = ((mul_22_25_n_788 & mul_22_25_n_746) | (mul_22_25_n_825 & (mul_22_25_n_788
    ^ mul_22_25_n_746)));
 assign mul_22_25_n_2009 = (mul_22_25_n_825 ^ (mul_22_25_n_788 ^ mul_22_25_n_746));
 assign mul_22_25_n_1992 = ((mul_22_25_n_992 & mul_22_25_n_956) | (mul_22_25_n_651 & (mul_22_25_n_992
    ^ mul_22_25_n_956)));
 assign mul_22_25_n_2010 = (mul_22_25_n_651 ^ (mul_22_25_n_992 ^ mul_22_25_n_956));
 assign mul_22_25_n_1991 = ((mul_22_25_n_760 & mul_22_25_n_718) | (mul_22_25_n_993 & (mul_22_25_n_760
    ^ mul_22_25_n_718)));
 assign mul_22_25_n_2008 = (mul_22_25_n_993 ^ (mul_22_25_n_760 ^ mul_22_25_n_718));
 assign mul_22_25_n_1986 = ((mul_22_25_n_1003 & mul_22_25_n_696) | (mul_22_25_n_1149 & (mul_22_25_n_1003
    ^ mul_22_25_n_696)));
 assign mul_22_25_n_2007 = (mul_22_25_n_1149 ^ (mul_22_25_n_1003 ^ mul_22_25_n_696));
 assign mul_22_25_n_1984 = ((mul_22_25_n_2014 & mul_22_25_n_2015) | (mul_22_25_n_2013 & (mul_22_25_n_2014
    ^ mul_22_25_n_2015)));
 assign mul_22_25_n_2003 = (mul_22_25_n_2013 ^ (mul_22_25_n_2014 ^ mul_22_25_n_2015));
 assign mul_22_25_n_1983 = ((mul_22_25_n_2011 & mul_22_25_n_2012) | (mul_22_25_n_2010 & (mul_22_25_n_2011
    ^ mul_22_25_n_2012)));
 assign mul_22_25_n_2001 = (mul_22_25_n_2010 ^ (mul_22_25_n_2011 ^ mul_22_25_n_2012));
 assign mul_22_25_n_1981 = ((mul_22_25_n_2008 & mul_22_25_n_2009) | (mul_22_25_n_2007 & (mul_22_25_n_2008
    ^ mul_22_25_n_2009)));
 assign mul_22_25_n_2002 = (mul_22_25_n_2007 ^ (mul_22_25_n_2008 ^ mul_22_25_n_2009));
 assign mul_22_25_n_1978 = ((mul_22_25_n_2005 & mul_22_25_n_2006) | (mul_22_25_n_2004 & (mul_22_25_n_2005
    ^ mul_22_25_n_2006)));
 assign mul_22_25_n_1999 = (mul_22_25_n_2004 ^ (mul_22_25_n_2005 ^ mul_22_25_n_2006));
 assign mul_22_25_n_1977 = ((mul_22_25_n_2002 & mul_22_25_n_2003) | (mul_22_25_n_2001 & (mul_22_25_n_2002
    ^ mul_22_25_n_2003)));
 assign mul_22_25_n_1997 = (mul_22_25_n_2001 ^ (mul_22_25_n_2002 ^ mul_22_25_n_2003));
 assign mul_22_25_n_1974 = ((mul_22_25_n_1999 & mul_22_25_n_2000) | (mul_22_25_n_1998 & (mul_22_25_n_1999
    ^ mul_22_25_n_2000)));
 assign mul_22_25_n_1995 = (mul_22_25_n_1998 ^ (mul_22_25_n_1999 ^ mul_22_25_n_2000));
 assign mul_22_25_n_2281 = ((n_72 & n_129) | (n_164 & (n_72 ^ n_129)));
 assign mul_22_25_n_2241 = (n_164 ^ (n_72 ^ n_129));
 assign mul_22_25_n_1972 = ((mul_22_25_n_706 & mul_22_25_n_1013) | (mul_22_25_n_1053 & (mul_22_25_n_706
    ^ mul_22_25_n_1013)));
 assign mul_22_25_n_1989 = (mul_22_25_n_1053 ^ (mul_22_25_n_706 ^ mul_22_25_n_1013));
 assign mul_22_25_n_1971 = ((mul_22_25_n_840 & mul_22_25_n_1107) | (mul_22_25_n_1047 & (mul_22_25_n_840
    ^ mul_22_25_n_1107)));
 assign mul_22_25_n_1987 = (mul_22_25_n_1047 ^ (mul_22_25_n_840 ^ mul_22_25_n_1107));
 assign mul_22_25_n_1969 = ((mul_22_25_n_783 & mul_22_25_n_682) | (mul_22_25_n_839 & (mul_22_25_n_783
    ^ mul_22_25_n_682)));
 assign mul_22_25_n_1988 = (mul_22_25_n_839 ^ (mul_22_25_n_783 ^ mul_22_25_n_682));
 assign mul_22_25_n_1970 = ((mul_22_25_n_1040 & mul_22_25_n_855) | (mul_22_25_n_1069 & (mul_22_25_n_1040
    ^ mul_22_25_n_855)));
 assign mul_22_25_n_1990 = (mul_22_25_n_1069 ^ (mul_22_25_n_1040 ^ mul_22_25_n_855));
 assign mul_22_25_n_1962 = ((mul_22_25_n_1176 & mul_22_25_n_1032) | (mul_22_25_n_1994 & (mul_22_25_n_1176
    ^ mul_22_25_n_1032)));
 assign mul_22_25_n_1985 = (mul_22_25_n_1994 ^ (mul_22_25_n_1176 ^ mul_22_25_n_1032));
 assign mul_22_25_n_1963 = ((mul_22_25_n_1992 & mul_22_25_n_1993) | (mul_22_25_n_1991 & (mul_22_25_n_1992
    ^ mul_22_25_n_1993)));
 assign mul_22_25_n_1982 = (mul_22_25_n_1991 ^ (mul_22_25_n_1992 ^ mul_22_25_n_1993));
 assign mul_22_25_n_1959 = ((mul_22_25_n_1989 & mul_22_25_n_1990) | (mul_22_25_n_1988 & (mul_22_25_n_1989
    ^ mul_22_25_n_1990)));
 assign mul_22_25_n_1980 = (mul_22_25_n_1988 ^ (mul_22_25_n_1989 ^ mul_22_25_n_1990));
 assign mul_22_25_n_1957 = ((mul_22_25_n_1986 & mul_22_25_n_1987) | (mul_22_25_n_1985 & (mul_22_25_n_1986
    ^ mul_22_25_n_1987)));
 assign mul_22_25_n_1979 = (mul_22_25_n_1985 ^ (mul_22_25_n_1986 ^ mul_22_25_n_1987));
 assign mul_22_25_n_1956 = ((mul_22_25_n_1983 & mul_22_25_n_1984) | (mul_22_25_n_1982 & (mul_22_25_n_1983
    ^ mul_22_25_n_1984)));
 assign mul_22_25_n_1976 = (mul_22_25_n_1982 ^ (mul_22_25_n_1983 ^ mul_22_25_n_1984));
 assign mul_22_25_n_1953 = ((mul_22_25_n_1980 & mul_22_25_n_1981) | (mul_22_25_n_1979 & (mul_22_25_n_1980
    ^ mul_22_25_n_1981)));
 assign mul_22_25_n_1975 = (mul_22_25_n_1979 ^ (mul_22_25_n_1980 ^ mul_22_25_n_1981));
 assign mul_22_25_n_1951 = ((mul_22_25_n_1977 & mul_22_25_n_1978) | (mul_22_25_n_1976 & (mul_22_25_n_1977
    ^ mul_22_25_n_1978)));
 assign mul_22_25_n_1973 = (mul_22_25_n_1976 ^ (mul_22_25_n_1977 ^ mul_22_25_n_1978));
 assign mul_22_25_n_2282 = ((n_165 & n_97) | (n_127 & (n_165 ^ n_97)));
 assign mul_22_25_n_2242 = (n_127 ^ (n_165 ^ n_97));
 assign mul_22_25_n_1948 = ((mul_22_25_n_900 & mul_22_25_n_636) | (mul_22_25_n_1012 & (mul_22_25_n_900
    ^ mul_22_25_n_636)));
 assign mul_22_25_n_1966 = (mul_22_25_n_1012 ^ (mul_22_25_n_900 ^ mul_22_25_n_636));
 assign mul_22_25_n_1947 = ((mul_22_25_n_742 & mul_22_25_n_965) | (mul_22_25_n_820 & (mul_22_25_n_742
    ^ mul_22_25_n_965)));
 assign mul_22_25_n_1968 = (mul_22_25_n_820 ^ (mul_22_25_n_742 ^ mul_22_25_n_965));
 assign mul_22_25_n_1949 = ((mul_22_25_n_980 & mul_22_25_n_989) | (mul_22_25_n_646 & (mul_22_25_n_980
    ^ mul_22_25_n_989)));
 assign mul_22_25_n_1965 = (mul_22_25_n_646 ^ (mul_22_25_n_980 ^ mul_22_25_n_989));
 assign mul_22_25_n_1946 = ((mul_22_25_n_1016 & mul_22_25_n_958) | (mul_22_25_n_743 & (mul_22_25_n_1016
    ^ mul_22_25_n_958)));
 assign mul_22_25_n_1964 = (mul_22_25_n_743 ^ (mul_22_25_n_1016 ^ mul_22_25_n_958));
 assign mul_22_25_n_1945 = ((mul_22_25_n_995 & mul_22_25_n_876) | (mul_22_25_n_994 & (mul_22_25_n_995
    ^ mul_22_25_n_876)));
 assign mul_22_25_n_1967 = (mul_22_25_n_994 ^ (mul_22_25_n_995 ^ mul_22_25_n_876));
 assign mul_22_25_n_1939 = ((mul_22_25_n_1972 & mul_22_25_n_1150) | (mul_22_25_n_1971 & (mul_22_25_n_1972
    ^ mul_22_25_n_1150)));
 assign mul_22_25_n_1961 = (mul_22_25_n_1971 ^ (mul_22_25_n_1972 ^ mul_22_25_n_1150));
 assign mul_22_25_n_1936 = ((mul_22_25_n_1969 & mul_22_25_n_1970) | (mul_22_25_n_1968 & (mul_22_25_n_1969
    ^ mul_22_25_n_1970)));
 assign mul_22_25_n_1960 = (mul_22_25_n_1968 ^ (mul_22_25_n_1969 ^ mul_22_25_n_1970));
 assign mul_22_25_n_1938 = ((mul_22_25_n_1966 & mul_22_25_n_1967) | (mul_22_25_n_1965 & (mul_22_25_n_1966
    ^ mul_22_25_n_1967)));
 assign mul_22_25_n_1958 = (mul_22_25_n_1965 ^ (mul_22_25_n_1966 ^ mul_22_25_n_1967));
 assign mul_22_25_n_1933 = ((mul_22_25_n_1963 & mul_22_25_n_1964) | (mul_22_25_n_1962 & (mul_22_25_n_1963
    ^ mul_22_25_n_1964)));
 assign mul_22_25_n_1955 = (mul_22_25_n_1962 ^ (mul_22_25_n_1963 ^ mul_22_25_n_1964));
 assign mul_22_25_n_1932 = ((mul_22_25_n_1960 & mul_22_25_n_1961) | (mul_22_25_n_1959 & (mul_22_25_n_1960
    ^ mul_22_25_n_1961)));
 assign mul_22_25_n_1954 = (mul_22_25_n_1959 ^ (mul_22_25_n_1960 ^ mul_22_25_n_1961));
 assign mul_22_25_n_1928 = ((mul_22_25_n_1957 & mul_22_25_n_1958) | (mul_22_25_n_1956 & (mul_22_25_n_1957
    ^ mul_22_25_n_1958)));
 assign mul_22_25_n_1952 = (mul_22_25_n_1956 ^ (mul_22_25_n_1957 ^ mul_22_25_n_1958));
 assign mul_22_25_n_1927 = ((mul_22_25_n_1954 & mul_22_25_n_1955) | (mul_22_25_n_1953 & (mul_22_25_n_1954
    ^ mul_22_25_n_1955)));
 assign mul_22_25_n_1950 = (mul_22_25_n_1953 ^ (mul_22_25_n_1954 ^ mul_22_25_n_1955));
 assign mul_22_25_n_2283 = ((n_128 & n_73) | (n_125 & (n_128 ^ n_73)));
 assign mul_22_25_n_2243 = (n_125 ^ (n_128 ^ n_73));
 assign mul_22_25_n_1925 = ((mul_22_25_n_863 & mul_22_25_n_978) | (mul_22_25_n_976 & (mul_22_25_n_863
    ^ mul_22_25_n_978)));
 assign mul_22_25_n_1944 = (mul_22_25_n_976 ^ (mul_22_25_n_863 ^ mul_22_25_n_978));
 assign mul_22_25_n_1924 = ((mul_22_25_n_961 & mul_22_25_n_709) | (mul_22_25_n_764 & (mul_22_25_n_961
    ^ mul_22_25_n_709)));
 assign mul_22_25_n_1942 = (mul_22_25_n_764 ^ (mul_22_25_n_961 ^ mul_22_25_n_709));
 assign mul_22_25_n_1923 = ((mul_22_25_n_968 & mul_22_25_n_1106) | (mul_22_25_n_765 & (mul_22_25_n_968
    ^ mul_22_25_n_1106)));
 assign mul_22_25_n_1941 = (mul_22_25_n_765 ^ (mul_22_25_n_968 ^ mul_22_25_n_1106));
 assign mul_22_25_n_1922 = ((mul_22_25_n_963 & mul_22_25_n_712) | (mul_22_25_n_974 & (mul_22_25_n_963
    ^ mul_22_25_n_712)));
 assign mul_22_25_n_1943 = (mul_22_25_n_974 ^ (mul_22_25_n_963 ^ mul_22_25_n_712));
 assign mul_22_25_n_1916 = ((mul_22_25_n_1070 & mul_22_25_n_999) | (mul_22_25_n_1165 & (mul_22_25_n_1070
    ^ mul_22_25_n_999)));
 assign mul_22_25_n_1940 = (mul_22_25_n_1165 ^ (mul_22_25_n_1070 ^ mul_22_25_n_999));
 assign mul_22_25_n_1914 = ((mul_22_25_n_1948 & mul_22_25_n_1949) | (mul_22_25_n_1947 & (mul_22_25_n_1948
    ^ mul_22_25_n_1949)));
 assign mul_22_25_n_1937 = (mul_22_25_n_1947 ^ (mul_22_25_n_1948 ^ mul_22_25_n_1949));
 assign mul_22_25_n_1911 = ((mul_22_25_n_1945 & mul_22_25_n_1946) | (mul_22_25_n_1944 & (mul_22_25_n_1945
    ^ mul_22_25_n_1946)));
 assign mul_22_25_n_1935 = (mul_22_25_n_1944 ^ (mul_22_25_n_1945 ^ mul_22_25_n_1946));
 assign mul_22_25_n_1913 = ((mul_22_25_n_1942 & mul_22_25_n_1943) | (mul_22_25_n_1941 & (mul_22_25_n_1942
    ^ mul_22_25_n_1943)));
 assign mul_22_25_n_1934 = (mul_22_25_n_1941 ^ (mul_22_25_n_1942 ^ mul_22_25_n_1943));
 assign mul_22_25_n_1907 = ((mul_22_25_n_1939 & mul_22_25_n_1940) | (mul_22_25_n_1938 & (mul_22_25_n_1939
    ^ mul_22_25_n_1940)));
 assign mul_22_25_n_1931 = (mul_22_25_n_1938 ^ (mul_22_25_n_1939 ^ mul_22_25_n_1940));
 assign mul_22_25_n_1908 = ((mul_22_25_n_1936 & mul_22_25_n_1937) | (mul_22_25_n_1935 & (mul_22_25_n_1936
    ^ mul_22_25_n_1937)));
 assign mul_22_25_n_1930 = (mul_22_25_n_1935 ^ (mul_22_25_n_1936 ^ mul_22_25_n_1937));
 assign mul_22_25_n_1904 = ((mul_22_25_n_1933 & mul_22_25_n_1934) | (mul_22_25_n_1932 & (mul_22_25_n_1933
    ^ mul_22_25_n_1934)));
 assign mul_22_25_n_1929 = (mul_22_25_n_1932 ^ (mul_22_25_n_1933 ^ mul_22_25_n_1934));
 assign mul_22_25_n_1901 = ((n_121 & n_110) | (n_69 & (n_121 ^ n_110)));
 assign mul_22_25_n_1926 = (n_69 ^ (n_121 ^ n_110));
 assign mul_22_25_n_2284 = ((n_126 & n_74) | (mul_22_25_n_1926 & (n_126 ^ n_74)));
 assign mul_22_25_n_2244 = (mul_22_25_n_1926 ^ (n_126 ^ n_74));
 assign mul_22_25_n_1900 = ((mul_22_25_n_652 & mul_22_25_n_633) | (mul_22_25_n_947 & (mul_22_25_n_652
    ^ mul_22_25_n_633)));
 assign mul_22_25_n_1921 = (mul_22_25_n_947 ^ (mul_22_25_n_652 ^ mul_22_25_n_633));
 assign mul_22_25_n_1899 = ((mul_22_25_n_945 & mul_22_25_n_874) | (mul_22_25_n_944 & (mul_22_25_n_945
    ^ mul_22_25_n_874)));
 assign mul_22_25_n_1917 = (mul_22_25_n_944 ^ (mul_22_25_n_945 ^ mul_22_25_n_874));
 assign mul_22_25_n_1898 = ((mul_22_25_n_1008 & mul_22_25_n_943) | (mul_22_25_n_941 & (mul_22_25_n_1008
    ^ mul_22_25_n_943)));
 assign mul_22_25_n_1918 = (mul_22_25_n_941 ^ (mul_22_25_n_1008 ^ mul_22_25_n_943));
 assign mul_22_25_n_1897 = ((mul_22_25_n_937 & mul_22_25_n_940) | (mul_22_25_n_936 & (mul_22_25_n_937
    ^ mul_22_25_n_940)));
 assign mul_22_25_n_1919 = (mul_22_25_n_936 ^ (mul_22_25_n_937 ^ mul_22_25_n_940));
 assign mul_22_25_n_1896 = ((mul_22_25_n_700 & mul_22_25_n_692) | (mul_22_25_n_931 & (mul_22_25_n_700
    ^ mul_22_25_n_692)));
 assign mul_22_25_n_1920 = (mul_22_25_n_931 ^ (mul_22_25_n_700 ^ mul_22_25_n_692));
 assign mul_22_25_n_1889 = ((mul_22_25_n_1160 & mul_22_25_n_929) | (mul_22_25_n_1925 & (mul_22_25_n_1160
    ^ mul_22_25_n_929)));
 assign mul_22_25_n_1915 = (mul_22_25_n_1925 ^ (mul_22_25_n_1160 ^ mul_22_25_n_929));
 assign mul_22_25_n_1890 = ((mul_22_25_n_1923 & mul_22_25_n_1924) | (mul_22_25_n_1922 & (mul_22_25_n_1923
    ^ mul_22_25_n_1924)));
 assign mul_22_25_n_1912 = (mul_22_25_n_1922 ^ (mul_22_25_n_1923 ^ mul_22_25_n_1924));
 assign mul_22_25_n_1886 = ((mul_22_25_n_1920 & mul_22_25_n_1921) | (mul_22_25_n_1919 & (mul_22_25_n_1920
    ^ mul_22_25_n_1921)));
 assign mul_22_25_n_1909 = (mul_22_25_n_1919 ^ (mul_22_25_n_1920 ^ mul_22_25_n_1921));
 assign mul_22_25_n_1885 = ((mul_22_25_n_1917 & mul_22_25_n_1918) | (mul_22_25_n_1916 & (mul_22_25_n_1917
    ^ mul_22_25_n_1918)));
 assign mul_22_25_n_1910 = (mul_22_25_n_1916 ^ (mul_22_25_n_1917 ^ mul_22_25_n_1918));
 assign mul_22_25_n_1882 = ((mul_22_25_n_1914 & mul_22_25_n_1915) | (mul_22_25_n_1913 & (mul_22_25_n_1914
    ^ mul_22_25_n_1915)));
 assign mul_22_25_n_1906 = (mul_22_25_n_1913 ^ (mul_22_25_n_1914 ^ mul_22_25_n_1915));
 assign mul_22_25_n_1881 = ((mul_22_25_n_1911 & mul_22_25_n_1912) | (mul_22_25_n_1910 & (mul_22_25_n_1911
    ^ mul_22_25_n_1912)));
 assign mul_22_25_n_1905 = (mul_22_25_n_1910 ^ (mul_22_25_n_1911 ^ mul_22_25_n_1912));
 assign mul_22_25_n_1878 = ((mul_22_25_n_1908 & mul_22_25_n_1909) | (mul_22_25_n_1907 & (mul_22_25_n_1908
    ^ mul_22_25_n_1909)));
 assign mul_22_25_n_1903 = (mul_22_25_n_1907 ^ (mul_22_25_n_1908 ^ mul_22_25_n_1909));
 assign mul_22_25_n_1875 = ((n_160 & n_106) | (n_70 & (n_160 ^ n_106)));
 assign mul_22_25_n_1902 = (n_70 ^ (n_160 ^ n_106));
 assign mul_22_25_n_2285 = ((mul_22_25_n_1902 & n_63) | (mul_22_25_n_1901 & (mul_22_25_n_1902 ^ n_63)));
 assign mul_22_25_n_2245 = (mul_22_25_n_1901 ^ (mul_22_25_n_1902 ^ n_63));
 assign mul_22_25_n_1874 = ((mul_22_25_n_1086 & mul_22_25_n_1110) | (mul_22_25_n_1071 & (mul_22_25_n_1086
    ^ mul_22_25_n_1110)));
 assign mul_22_25_n_1894 = (mul_22_25_n_1071 ^ (mul_22_25_n_1086 ^ mul_22_25_n_1110));
 assign mul_22_25_n_1873 = ((mul_22_25_n_1095 & mul_22_25_n_1093) | (mul_22_25_n_1096 & (mul_22_25_n_1095
    ^ mul_22_25_n_1093)));
 assign mul_22_25_n_1893 = (mul_22_25_n_1096 ^ (mul_22_25_n_1095 ^ mul_22_25_n_1093));
 assign mul_22_25_n_1872 = ((mul_22_25_n_1098 & mul_22_25_n_1097) | (mul_22_25_n_1100 & (mul_22_25_n_1098
    ^ mul_22_25_n_1097)));
 assign mul_22_25_n_1892 = (mul_22_25_n_1100 ^ (mul_22_25_n_1098 ^ mul_22_25_n_1097));
 assign mul_22_25_n_1871 = ((mul_22_25_n_1104 & mul_22_25_n_1034) | (mul_22_25_n_1051 & (mul_22_25_n_1104
    ^ mul_22_25_n_1034)));
 assign mul_22_25_n_1891 = (mul_22_25_n_1051 ^ (mul_22_25_n_1104 ^ mul_22_25_n_1034));
 assign mul_22_25_n_1870 = ((mul_22_25_n_710 & mul_22_25_n_1111) | (mul_22_25_n_1112 & (mul_22_25_n_710
    ^ mul_22_25_n_1111)));
 assign mul_22_25_n_1895 = (mul_22_25_n_1112 ^ (mul_22_25_n_710 ^ mul_22_25_n_1111));
 assign mul_22_25_n_1863 = ((mul_22_25_n_1900 & mul_22_25_n_1177) | (mul_22_25_n_1899 & (mul_22_25_n_1900
    ^ mul_22_25_n_1177)));
 assign mul_22_25_n_1887 = (mul_22_25_n_1899 ^ (mul_22_25_n_1900 ^ mul_22_25_n_1177));
 assign mul_22_25_n_1864 = ((mul_22_25_n_1897 & mul_22_25_n_1898) | (mul_22_25_n_1896 & (mul_22_25_n_1897
    ^ mul_22_25_n_1898)));
 assign mul_22_25_n_1888 = (mul_22_25_n_1896 ^ (mul_22_25_n_1897 ^ mul_22_25_n_1898));
 assign mul_22_25_n_1862 = ((mul_22_25_n_1894 & mul_22_25_n_1895) | (mul_22_25_n_1893 & (mul_22_25_n_1894
    ^ mul_22_25_n_1895)));
 assign mul_22_25_n_1884 = (mul_22_25_n_1893 ^ (mul_22_25_n_1894 ^ mul_22_25_n_1895));
 assign mul_22_25_n_1858 = ((mul_22_25_n_1891 & mul_22_25_n_1892) | (mul_22_25_n_1890 & (mul_22_25_n_1891
    ^ mul_22_25_n_1892)));
 assign mul_22_25_n_1883 = (mul_22_25_n_1890 ^ (mul_22_25_n_1891 ^ mul_22_25_n_1892));
 assign mul_22_25_n_1856 = ((mul_22_25_n_1888 & mul_22_25_n_1889) | (mul_22_25_n_1887 & (mul_22_25_n_1888
    ^ mul_22_25_n_1889)));
 assign mul_22_25_n_1880 = (mul_22_25_n_1887 ^ (mul_22_25_n_1888 ^ mul_22_25_n_1889));
 assign mul_22_25_n_1855 = ((mul_22_25_n_1885 & mul_22_25_n_1886) | (mul_22_25_n_1884 & (mul_22_25_n_1885
    ^ mul_22_25_n_1886)));
 assign mul_22_25_n_1879 = (mul_22_25_n_1884 ^ (mul_22_25_n_1885 ^ mul_22_25_n_1886));
 assign mul_22_25_n_1851 = ((mul_22_25_n_1882 & mul_22_25_n_1883) | (mul_22_25_n_1881 & (mul_22_25_n_1882
    ^ mul_22_25_n_1883)));
 assign mul_22_25_n_1877 = (mul_22_25_n_1881 ^ (mul_22_25_n_1882 ^ mul_22_25_n_1883));
 assign mul_22_25_n_1850 = ((n_77 & n_100) | (n_64 & (n_77 ^ n_100)));
 assign mul_22_25_n_1876 = (n_64 ^ (n_77 ^ n_100));
 assign mul_22_25_n_2286 = ((mul_22_25_n_1876 & n_158) | (mul_22_25_n_1875 & (mul_22_25_n_1876 ^ n_158)));
 assign mul_22_25_n_2246 = (mul_22_25_n_1875 ^ (mul_22_25_n_1876 ^ n_158));
 assign mul_22_25_n_1848 = ((mul_22_25_n_894 & mul_22_25_n_895) | (mul_22_25_n_893 & (mul_22_25_n_894
    ^ mul_22_25_n_895)));
 assign mul_22_25_n_1866 = (mul_22_25_n_893 ^ (mul_22_25_n_894 ^ mul_22_25_n_895));
 assign mul_22_25_n_1847 = ((mul_22_25_n_892 & mul_22_25_n_960) | (mul_22_25_n_891 & (mul_22_25_n_892
    ^ mul_22_25_n_960)));
 assign mul_22_25_n_1869 = (mul_22_25_n_891 ^ (mul_22_25_n_892 ^ mul_22_25_n_960));
 assign mul_22_25_n_1846 = ((mul_22_25_n_887 & mul_22_25_n_889) | (mul_22_25_n_885 & (mul_22_25_n_887
    ^ mul_22_25_n_889)));
 assign mul_22_25_n_1868 = (mul_22_25_n_885 ^ (mul_22_25_n_887 ^ mul_22_25_n_889));
 assign mul_22_25_n_1845 = ((mul_22_25_n_881 & mul_22_25_n_882) | (mul_22_25_n_880 & (mul_22_25_n_881
    ^ mul_22_25_n_882)));
 assign mul_22_25_n_1867 = (mul_22_25_n_880 ^ (mul_22_25_n_881 ^ mul_22_25_n_882));
 assign mul_22_25_n_1839 = ((mul_22_25_n_877 & mul_22_25_n_878) | (mul_22_25_n_1144 & (mul_22_25_n_877
    ^ mul_22_25_n_878)));
 assign mul_22_25_n_1865 = (mul_22_25_n_1144 ^ (mul_22_25_n_877 ^ mul_22_25_n_878));
 assign mul_22_25_n_1838 = ((mul_22_25_n_1873 & mul_22_25_n_1874) | (mul_22_25_n_1872 & (mul_22_25_n_1873
    ^ mul_22_25_n_1874)));
 assign mul_22_25_n_1860 = (mul_22_25_n_1872 ^ (mul_22_25_n_1873 ^ mul_22_25_n_1874));
 assign mul_22_25_n_1837 = ((mul_22_25_n_1870 & mul_22_25_n_1871) | (mul_22_25_n_1173 & (mul_22_25_n_1870
    ^ mul_22_25_n_1871)));
 assign mul_22_25_n_1861 = (mul_22_25_n_1173 ^ (mul_22_25_n_1870 ^ mul_22_25_n_1871));
 assign mul_22_25_n_1834 = ((mul_22_25_n_1868 & mul_22_25_n_1869) | (mul_22_25_n_1867 & (mul_22_25_n_1868
    ^ mul_22_25_n_1869)));
 assign mul_22_25_n_1859 = (mul_22_25_n_1867 ^ (mul_22_25_n_1868 ^ mul_22_25_n_1869));
 assign mul_22_25_n_1831 = ((mul_22_25_n_1865 & mul_22_25_n_1866) | (mul_22_25_n_1864 & (mul_22_25_n_1865
    ^ mul_22_25_n_1866)));
 assign mul_22_25_n_1857 = (mul_22_25_n_1864 ^ (mul_22_25_n_1865 ^ mul_22_25_n_1866));
 assign mul_22_25_n_1830 = ((mul_22_25_n_1862 & mul_22_25_n_1863) | (mul_22_25_n_1861 & (mul_22_25_n_1862
    ^ mul_22_25_n_1863)));
 assign mul_22_25_n_1854 = (mul_22_25_n_1861 ^ (mul_22_25_n_1862 ^ mul_22_25_n_1863));
 assign mul_22_25_n_1827 = ((mul_22_25_n_1859 & mul_22_25_n_1860) | (mul_22_25_n_1858 & (mul_22_25_n_1859
    ^ mul_22_25_n_1860)));
 assign mul_22_25_n_1853 = (mul_22_25_n_1858 ^ (mul_22_25_n_1859 ^ mul_22_25_n_1860));
 assign mul_22_25_n_1826 = ((mul_22_25_n_1856 & mul_22_25_n_1857) | (mul_22_25_n_1855 & (mul_22_25_n_1856
    ^ mul_22_25_n_1857)));
 assign mul_22_25_n_1852 = (mul_22_25_n_1855 ^ (mul_22_25_n_1856 ^ mul_22_25_n_1857));
 assign mul_22_25_n_1823 = ((n_162 & n_68) | (n_98 & (n_162 ^ n_68)));
 assign mul_22_25_n_1849 = (n_98 ^ (n_162 ^ n_68));
 assign mul_22_25_n_2287 = ((mul_22_25_n_1850 & n_159) | (mul_22_25_n_1849 & (mul_22_25_n_1850 ^ n_159)));
 assign mul_22_25_n_2247 = (mul_22_25_n_1849 ^ (mul_22_25_n_1850 ^ n_159));
 assign mul_22_25_n_1822 = ((mul_22_25_n_857 & mul_22_25_n_883) | (mul_22_25_n_856 & (mul_22_25_n_857
    ^ mul_22_25_n_883)));
 assign mul_22_25_n_1844 = (mul_22_25_n_856 ^ (mul_22_25_n_857 ^ mul_22_25_n_883));
 assign mul_22_25_n_1821 = ((mul_22_25_n_853 & mul_22_25_n_998) | (mul_22_25_n_852 & (mul_22_25_n_853
    ^ mul_22_25_n_998)));
 assign mul_22_25_n_1842 = (mul_22_25_n_852 ^ (mul_22_25_n_853 ^ mul_22_25_n_998));
 assign mul_22_25_n_1820 = ((mul_22_25_n_850 & mul_22_25_n_851) | (mul_22_25_n_966 & (mul_22_25_n_850
    ^ mul_22_25_n_851)));
 assign mul_22_25_n_1841 = (mul_22_25_n_966 ^ (mul_22_25_n_850 ^ mul_22_25_n_851));
 assign mul_22_25_n_1819 = ((mul_22_25_n_848 & mul_22_25_n_1048) | (mul_22_25_n_847 & (mul_22_25_n_848
    ^ mul_22_25_n_1048)));
 assign mul_22_25_n_1843 = (mul_22_25_n_847 ^ (mul_22_25_n_848 ^ mul_22_25_n_1048));
 assign mul_22_25_n_1813 = ((mul_22_25_n_842 & mul_22_25_n_1022) | (mul_22_25_n_1139 & (mul_22_25_n_842
    ^ mul_22_25_n_1022)));
 assign mul_22_25_n_1840 = (mul_22_25_n_1139 ^ (mul_22_25_n_842 ^ mul_22_25_n_1022));
 assign mul_22_25_n_1812 = ((mul_22_25_n_1848 & mul_22_25_n_1152) | (mul_22_25_n_1847 & (mul_22_25_n_1848
    ^ mul_22_25_n_1152)));
 assign mul_22_25_n_1836 = (mul_22_25_n_1847 ^ (mul_22_25_n_1848 ^ mul_22_25_n_1152));
 assign mul_22_25_n_1809 = ((mul_22_25_n_1845 & mul_22_25_n_1846) | (mul_22_25_n_1844 & (mul_22_25_n_1845
    ^ mul_22_25_n_1846)));
 assign mul_22_25_n_1835 = (mul_22_25_n_1844 ^ (mul_22_25_n_1845 ^ mul_22_25_n_1846));
 assign mul_22_25_n_1808 = ((mul_22_25_n_1842 & mul_22_25_n_1843) | (mul_22_25_n_1841 & (mul_22_25_n_1842
    ^ mul_22_25_n_1843)));
 assign mul_22_25_n_1833 = (mul_22_25_n_1841 ^ (mul_22_25_n_1842 ^ mul_22_25_n_1843));
 assign mul_22_25_n_1805 = ((mul_22_25_n_1839 & mul_22_25_n_1840) | (mul_22_25_n_1838 & (mul_22_25_n_1839
    ^ mul_22_25_n_1840)));
 assign mul_22_25_n_1832 = (mul_22_25_n_1838 ^ (mul_22_25_n_1839 ^ mul_22_25_n_1840));
 assign mul_22_25_n_1804 = ((mul_22_25_n_1836 & mul_22_25_n_1837) | (mul_22_25_n_1835 & (mul_22_25_n_1836
    ^ mul_22_25_n_1837)));
 assign mul_22_25_n_1829 = (mul_22_25_n_1835 ^ (mul_22_25_n_1836 ^ mul_22_25_n_1837));
 assign mul_22_25_n_1801 = ((mul_22_25_n_1833 & mul_22_25_n_1834) | (mul_22_25_n_1832 & (mul_22_25_n_1833
    ^ mul_22_25_n_1834)));
 assign mul_22_25_n_1828 = (mul_22_25_n_1832 ^ (mul_22_25_n_1833 ^ mul_22_25_n_1834));
 assign mul_22_25_n_1800 = ((mul_22_25_n_1830 & mul_22_25_n_1831) | (mul_22_25_n_1829 & (mul_22_25_n_1830
    ^ mul_22_25_n_1831)));
 assign mul_22_25_n_1825 = (mul_22_25_n_1829 ^ (mul_22_25_n_1830 ^ mul_22_25_n_1831));
 assign mul_22_25_n_1797 = ((n_163 & n_75) | (n_99 & (n_163 ^ n_75)));
 assign mul_22_25_n_1824 = (n_99 ^ (n_163 ^ n_75));
 assign mul_22_25_n_2288 = ((mul_22_25_n_1824 & n_117) | (mul_22_25_n_1823 & (mul_22_25_n_1824 ^ n_117)));
 assign mul_22_25_n_2248 = (mul_22_25_n_1823 ^ (mul_22_25_n_1824 ^ n_117));
 assign mul_22_25_n_1795 = ((mul_22_25_n_824 & mul_22_25_n_1085) | (mul_22_25_n_822 & (mul_22_25_n_824
    ^ mul_22_25_n_1085)));
 assign mul_22_25_n_1816 = (mul_22_25_n_822 ^ (mul_22_25_n_824 ^ mul_22_25_n_1085));
 assign mul_22_25_n_1794 = ((mul_22_25_n_819 & mul_22_25_n_821) | (mul_22_25_n_1029 & (mul_22_25_n_819
    ^ mul_22_25_n_821)));
 assign mul_22_25_n_1818 = (mul_22_25_n_1029 ^ (mul_22_25_n_819 ^ mul_22_25_n_821));
 assign mul_22_25_n_1793 = ((mul_22_25_n_690 & mul_22_25_n_715) | (mul_22_25_n_817 & (mul_22_25_n_690
    ^ mul_22_25_n_715)));
 assign mul_22_25_n_1814 = (mul_22_25_n_817 ^ (mul_22_25_n_690 ^ mul_22_25_n_715));
 assign mul_22_25_n_1796 = ((mul_22_25_n_811 & mul_22_25_n_719) | (mul_22_25_n_724 & (mul_22_25_n_811
    ^ mul_22_25_n_719)));
 assign mul_22_25_n_1815 = (mul_22_25_n_724 ^ (mul_22_25_n_811 ^ mul_22_25_n_719));
 assign mul_22_25_n_1792 = ((mul_22_25_n_808 & mul_22_25_n_809) | (mul_22_25_n_807 & (mul_22_25_n_808
    ^ mul_22_25_n_809)));
 assign mul_22_25_n_1817 = (mul_22_25_n_807 ^ (mul_22_25_n_808 ^ mul_22_25_n_809));
 assign mul_22_25_n_1786 = ((mul_22_25_n_1822 & mul_22_25_n_1140) | (mul_22_25_n_1821 & (mul_22_25_n_1822
    ^ mul_22_25_n_1140)));
 assign mul_22_25_n_1811 = (mul_22_25_n_1821 ^ (mul_22_25_n_1822 ^ mul_22_25_n_1140));
 assign mul_22_25_n_1784 = ((mul_22_25_n_1819 & mul_22_25_n_1820) | (mul_22_25_n_1818 & (mul_22_25_n_1819
    ^ mul_22_25_n_1820)));
 assign mul_22_25_n_1810 = (mul_22_25_n_1818 ^ (mul_22_25_n_1819 ^ mul_22_25_n_1820));
 assign mul_22_25_n_1783 = ((mul_22_25_n_1816 & mul_22_25_n_1817) | (mul_22_25_n_1815 & (mul_22_25_n_1816
    ^ mul_22_25_n_1817)));
 assign mul_22_25_n_1807 = (mul_22_25_n_1815 ^ (mul_22_25_n_1816 ^ mul_22_25_n_1817));
 assign mul_22_25_n_1781 = ((mul_22_25_n_1813 & mul_22_25_n_1814) | (mul_22_25_n_1812 & (mul_22_25_n_1813
    ^ mul_22_25_n_1814)));
 assign mul_22_25_n_1806 = (mul_22_25_n_1812 ^ (mul_22_25_n_1813 ^ mul_22_25_n_1814));
 assign mul_22_25_n_1779 = ((mul_22_25_n_1810 & mul_22_25_n_1811) | (mul_22_25_n_1809 & (mul_22_25_n_1810
    ^ mul_22_25_n_1811)));
 assign mul_22_25_n_1803 = (mul_22_25_n_1809 ^ (mul_22_25_n_1810 ^ mul_22_25_n_1811));
 assign mul_22_25_n_1776 = ((mul_22_25_n_1807 & mul_22_25_n_1808) | (mul_22_25_n_1806 & (mul_22_25_n_1807
    ^ mul_22_25_n_1808)));
 assign mul_22_25_n_1802 = (mul_22_25_n_1806 ^ (mul_22_25_n_1807 ^ mul_22_25_n_1808));
 assign mul_22_25_n_1774 = ((mul_22_25_n_1804 & mul_22_25_n_1805) | (mul_22_25_n_1803 & (mul_22_25_n_1804
    ^ mul_22_25_n_1805)));
 assign mul_22_25_n_1799 = (mul_22_25_n_1803 ^ (mul_22_25_n_1804 ^ mul_22_25_n_1805));
 assign mul_22_25_n_1772 = ((n_76 & n_119) | (n_118 & (n_76 ^ n_119)));
 assign mul_22_25_n_1798 = (n_118 ^ (n_76 ^ n_119));
 assign mul_22_25_n_2289 = ((mul_22_25_n_1798 & n_168) | (mul_22_25_n_1797 & (mul_22_25_n_1798 ^ n_168)));
 assign mul_22_25_n_2249 = (mul_22_25_n_1797 ^ (mul_22_25_n_1798 ^ n_168));
 assign mul_22_25_n_1771 = ((mul_22_25_n_802 & mul_22_25_n_973) | (mul_22_25_n_800 & (mul_22_25_n_802
    ^ mul_22_25_n_973)));
 assign mul_22_25_n_1790 = (mul_22_25_n_800 ^ (mul_22_25_n_802 ^ mul_22_25_n_973));
 assign mul_22_25_n_1770 = ((mul_22_25_n_1023 & mul_22_25_n_1056) | (mul_22_25_n_1028 & (mul_22_25_n_1023
    ^ mul_22_25_n_1056)));
 assign mul_22_25_n_1788 = (mul_22_25_n_1028 ^ (mul_22_25_n_1023 ^ mul_22_25_n_1056));
 assign mul_22_25_n_1769 = ((mul_22_25_n_797 & mul_22_25_n_1084) | (mul_22_25_n_796 & (mul_22_25_n_797
    ^ mul_22_25_n_1084)));
 assign mul_22_25_n_1789 = (mul_22_25_n_796 ^ (mul_22_25_n_797 ^ mul_22_25_n_1084));
 assign mul_22_25_n_1768 = ((mul_22_25_n_1054 & mul_22_25_n_767) | (mul_22_25_n_836 & (mul_22_25_n_1054
    ^ mul_22_25_n_767)));
 assign mul_22_25_n_1791 = (mul_22_25_n_836 ^ (mul_22_25_n_1054 ^ mul_22_25_n_767));
 assign mul_22_25_n_1762 = ((mul_22_25_n_913 & mul_22_25_n_794) | (mul_22_25_n_1796 & (mul_22_25_n_913
    ^ mul_22_25_n_794)));
 assign mul_22_25_n_1787 = (mul_22_25_n_1796 ^ (mul_22_25_n_913 ^ mul_22_25_n_794));
 assign mul_22_25_n_1761 = ((mul_22_25_n_1794 & mul_22_25_n_1795) | (mul_22_25_n_1793 & (mul_22_25_n_1794
    ^ mul_22_25_n_1795)));
 assign mul_22_25_n_1785 = (mul_22_25_n_1793 ^ (mul_22_25_n_1794 ^ mul_22_25_n_1795));
 assign mul_22_25_n_1759 = ((mul_22_25_n_1791 & mul_22_25_n_1792) | (mul_22_25_n_1790 & (mul_22_25_n_1791
    ^ mul_22_25_n_1792)));
 assign mul_22_25_n_1782 = (mul_22_25_n_1790 ^ (mul_22_25_n_1791 ^ mul_22_25_n_1792));
 assign mul_22_25_n_1756 = ((mul_22_25_n_1788 & mul_22_25_n_1789) | (mul_22_25_n_1787 & (mul_22_25_n_1788
    ^ mul_22_25_n_1789)));
 assign mul_22_25_n_1780 = (mul_22_25_n_1787 ^ (mul_22_25_n_1788 ^ mul_22_25_n_1789));
 assign mul_22_25_n_1754 = ((mul_22_25_n_1785 & mul_22_25_n_1786) | (mul_22_25_n_1784 & (mul_22_25_n_1785
    ^ mul_22_25_n_1786)));
 assign mul_22_25_n_1778 = (mul_22_25_n_1784 ^ (mul_22_25_n_1785 ^ mul_22_25_n_1786));
 assign mul_22_25_n_1753 = ((mul_22_25_n_1782 & mul_22_25_n_1783) | (mul_22_25_n_1781 & (mul_22_25_n_1782
    ^ mul_22_25_n_1783)));
 assign mul_22_25_n_1777 = (mul_22_25_n_1781 ^ (mul_22_25_n_1782 ^ mul_22_25_n_1783));
 assign mul_22_25_n_1750 = ((mul_22_25_n_1779 & mul_22_25_n_1780) | (mul_22_25_n_1778 & (mul_22_25_n_1779
    ^ mul_22_25_n_1780)));
 assign mul_22_25_n_1775 = (mul_22_25_n_1778 ^ (mul_22_25_n_1779 ^ mul_22_25_n_1780));
 assign mul_22_25_n_1748 = ((n_120 & n_102) | (n_140 & (n_120 ^ n_102)));
 assign mul_22_25_n_1773 = (n_140 ^ (n_120 ^ n_102));
 assign mul_22_25_n_2290 = ((mul_22_25_n_1773 & n_169) | (mul_22_25_n_1772 & (mul_22_25_n_1773 ^ n_169)));
 assign mul_22_25_n_2250 = (mul_22_25_n_1772 ^ (mul_22_25_n_1773 ^ n_169));
 assign mul_22_25_n_1744 = ((mul_22_25_n_781 & mul_22_25_n_1083) | (mul_22_25_n_933 & (mul_22_25_n_781
    ^ mul_22_25_n_1083)));
 assign mul_22_25_n_1766 = (mul_22_25_n_933 ^ (mul_22_25_n_781 ^ mul_22_25_n_1083));
 assign mul_22_25_n_1747 = ((mul_22_25_n_777 & mul_22_25_n_778) | (mul_22_25_n_948 & (mul_22_25_n_777
    ^ mul_22_25_n_778)));
 assign mul_22_25_n_1767 = (mul_22_25_n_948 ^ (mul_22_25_n_777 ^ mul_22_25_n_778));
 assign mul_22_25_n_1746 = ((mul_22_25_n_775 & mul_22_25_n_1045) | (mul_22_25_n_1108 & (mul_22_25_n_775
    ^ mul_22_25_n_1045)));
 assign mul_22_25_n_1764 = (mul_22_25_n_1108 ^ (mul_22_25_n_775 ^ mul_22_25_n_1045));
 assign mul_22_25_n_1745 = ((mul_22_25_n_770 & mul_22_25_n_772) | (mul_22_25_n_769 & (mul_22_25_n_770
    ^ mul_22_25_n_772)));
 assign mul_22_25_n_1765 = (mul_22_25_n_769 ^ (mul_22_25_n_770 ^ mul_22_25_n_772));
 assign mul_22_25_n_1739 = ((mul_22_25_n_698 & mul_22_25_n_834) | (mul_22_25_n_912 & (mul_22_25_n_698
    ^ mul_22_25_n_834)));
 assign mul_22_25_n_1763 = (mul_22_25_n_912 ^ (mul_22_25_n_698 ^ mul_22_25_n_834));
 assign mul_22_25_n_1738 = ((mul_22_25_n_1770 & mul_22_25_n_1771) | (mul_22_25_n_1769 & (mul_22_25_n_1770
    ^ mul_22_25_n_1771)));
 assign mul_22_25_n_1760 = (mul_22_25_n_1769 ^ (mul_22_25_n_1770 ^ mul_22_25_n_1771));
 assign mul_22_25_n_1735 = ((mul_22_25_n_1767 & mul_22_25_n_1768) | (mul_22_25_n_1766 & (mul_22_25_n_1767
    ^ mul_22_25_n_1768)));
 assign mul_22_25_n_1758 = (mul_22_25_n_1766 ^ (mul_22_25_n_1767 ^ mul_22_25_n_1768));
 assign mul_22_25_n_1734 = ((mul_22_25_n_1764 & mul_22_25_n_1765) | (mul_22_25_n_1763 & (mul_22_25_n_1764
    ^ mul_22_25_n_1765)));
 assign mul_22_25_n_1757 = (mul_22_25_n_1763 ^ (mul_22_25_n_1764 ^ mul_22_25_n_1765));
 assign mul_22_25_n_1732 = ((mul_22_25_n_1761 & mul_22_25_n_1762) | (mul_22_25_n_1760 & (mul_22_25_n_1761
    ^ mul_22_25_n_1762)));
 assign mul_22_25_n_1755 = (mul_22_25_n_1760 ^ (mul_22_25_n_1761 ^ mul_22_25_n_1762));
 assign mul_22_25_n_1729 = ((mul_22_25_n_1758 & mul_22_25_n_1759) | (mul_22_25_n_1757 & (mul_22_25_n_1758
    ^ mul_22_25_n_1759)));
 assign mul_22_25_n_1752 = (mul_22_25_n_1757 ^ (mul_22_25_n_1758 ^ mul_22_25_n_1759));
 assign mul_22_25_n_1728 = ((mul_22_25_n_1755 & mul_22_25_n_1756) | (mul_22_25_n_1754 & (mul_22_25_n_1755
    ^ mul_22_25_n_1756)));
 assign mul_22_25_n_1751 = (mul_22_25_n_1754 ^ (mul_22_25_n_1755 ^ mul_22_25_n_1756));
 assign mul_22_25_n_1725 = ((n_48 & n_103) | (n_146 & (n_48 ^ n_103)));
 assign mul_22_25_n_1749 = (n_146 ^ (n_48 ^ n_103));
 assign mul_22_25_n_2291 = ((mul_22_25_n_1749 & n_141) | (mul_22_25_n_1748 & (mul_22_25_n_1749 ^ n_141)));
 assign mul_22_25_n_2251 = (mul_22_25_n_1748 ^ (mul_22_25_n_1749 ^ n_141));
 assign mul_22_25_n_1721 = ((mul_22_25_n_986 & mul_22_25_n_762) | (mul_22_25_n_1004 & (mul_22_25_n_986
    ^ mul_22_25_n_762)));
 assign mul_22_25_n_1742 = (mul_22_25_n_1004 ^ (mul_22_25_n_986 ^ mul_22_25_n_762));
 assign mul_22_25_n_1724 = ((mul_22_25_n_761 & mul_22_25_n_983) | (mul_22_25_n_716 & (mul_22_25_n_761
    ^ mul_22_25_n_983)));
 assign mul_22_25_n_1740 = (mul_22_25_n_716 ^ (mul_22_25_n_761 ^ mul_22_25_n_983));
 assign mul_22_25_n_1723 = ((mul_22_25_n_727 & mul_22_25_n_1079) | (mul_22_25_n_757 & (mul_22_25_n_727
    ^ mul_22_25_n_1079)));
 assign mul_22_25_n_1741 = (mul_22_25_n_757 ^ (mul_22_25_n_727 ^ mul_22_25_n_1079));
 assign mul_22_25_n_1722 = ((mul_22_25_n_756 & mul_22_25_n_759) | (mul_22_25_n_789 & (mul_22_25_n_756
    ^ mul_22_25_n_759)));
 assign mul_22_25_n_1743 = (mul_22_25_n_789 ^ (mul_22_25_n_756 ^ mul_22_25_n_759));
 assign mul_22_25_n_1715 = ((mul_22_25_n_1747 & mul_22_25_n_916) | (mul_22_25_n_1746 & (mul_22_25_n_1747
    ^ mul_22_25_n_916)));
 assign mul_22_25_n_1737 = (mul_22_25_n_1746 ^ (mul_22_25_n_1747 ^ mul_22_25_n_916));
 assign mul_22_25_n_1713 = ((mul_22_25_n_1744 & mul_22_25_n_1745) | (mul_22_25_n_1743 & (mul_22_25_n_1744
    ^ mul_22_25_n_1745)));
 assign mul_22_25_n_1736 = (mul_22_25_n_1743 ^ (mul_22_25_n_1744 ^ mul_22_25_n_1745));
 assign mul_22_25_n_1712 = ((mul_22_25_n_1741 & mul_22_25_n_1742) | (mul_22_25_n_1740 & (mul_22_25_n_1741
    ^ mul_22_25_n_1742)));
 assign mul_22_25_n_1733 = (mul_22_25_n_1740 ^ (mul_22_25_n_1741 ^ mul_22_25_n_1742));
 assign mul_22_25_n_1710 = ((mul_22_25_n_1738 & mul_22_25_n_1739) | (mul_22_25_n_1737 & (mul_22_25_n_1738
    ^ mul_22_25_n_1739)));
 assign mul_22_25_n_1731 = (mul_22_25_n_1737 ^ (mul_22_25_n_1738 ^ mul_22_25_n_1739));
 assign mul_22_25_n_1708 = ((mul_22_25_n_1735 & mul_22_25_n_1736) | (mul_22_25_n_1734 & (mul_22_25_n_1735
    ^ mul_22_25_n_1736)));
 assign mul_22_25_n_1730 = (mul_22_25_n_1734 ^ (mul_22_25_n_1735 ^ mul_22_25_n_1736));
 assign mul_22_25_n_1706 = ((mul_22_25_n_1732 & mul_22_25_n_1733) | (mul_22_25_n_1731 & (mul_22_25_n_1732
    ^ mul_22_25_n_1733)));
 assign mul_22_25_n_1727 = (mul_22_25_n_1731 ^ (mul_22_25_n_1732 ^ mul_22_25_n_1733));
 assign mul_22_25_n_1703 = ((n_49 & n_172) | (n_147 & (n_49 ^ n_172)));
 assign mul_22_25_n_1726 = (n_147 ^ (n_49 ^ n_172));
 assign mul_22_25_n_2292 = ((mul_22_25_n_1726 & n_104) | (mul_22_25_n_1725 & (mul_22_25_n_1726 ^ n_104)));
 assign mul_22_25_n_2252 = (mul_22_25_n_1725 ^ (mul_22_25_n_1726 ^ n_104));
 assign mul_22_25_n_1700 = ((mul_22_25_n_741 & mul_22_25_n_1082) | (mul_22_25_n_1039 & (mul_22_25_n_741
    ^ mul_22_25_n_1082)));
 assign mul_22_25_n_1720 = (mul_22_25_n_1039 ^ (mul_22_25_n_741 ^ mul_22_25_n_1082));
 assign mul_22_25_n_1699 = ((mul_22_25_n_737 & mul_22_25_n_739) | (mul_22_25_n_736 & (mul_22_25_n_737
    ^ mul_22_25_n_739)));
 assign mul_22_25_n_1718 = (mul_22_25_n_736 ^ (mul_22_25_n_737 ^ mul_22_25_n_739));
 assign mul_22_25_n_1702 = ((mul_22_25_n_732 & mul_22_25_n_734) | (mul_22_25_n_731 & (mul_22_25_n_732
    ^ mul_22_25_n_734)));
 assign mul_22_25_n_1719 = (mul_22_25_n_731 ^ (mul_22_25_n_732 ^ mul_22_25_n_734));
 assign mul_22_25_n_1701 = ((mul_22_25_n_730 & mul_22_25_n_1102) | (mul_22_25_n_955 & (mul_22_25_n_730
    ^ mul_22_25_n_1102)));
 assign mul_22_25_n_1717 = (mul_22_25_n_955 ^ (mul_22_25_n_730 ^ mul_22_25_n_1102));
 assign mul_22_25_n_1693 = ((mul_22_25_n_915 & mul_22_25_n_728) | (mul_22_25_n_1724 & (mul_22_25_n_915
    ^ mul_22_25_n_728)));
 assign mul_22_25_n_1716 = (mul_22_25_n_1724 ^ (mul_22_25_n_915 ^ mul_22_25_n_728));
 assign mul_22_25_n_1694 = ((mul_22_25_n_1722 & mul_22_25_n_1723) | (mul_22_25_n_1721 & (mul_22_25_n_1722
    ^ mul_22_25_n_1723)));
 assign mul_22_25_n_1714 = (mul_22_25_n_1721 ^ (mul_22_25_n_1722 ^ mul_22_25_n_1723));
 assign mul_22_25_n_1691 = ((mul_22_25_n_1719 & mul_22_25_n_1720) | (mul_22_25_n_1718 & (mul_22_25_n_1719
    ^ mul_22_25_n_1720)));
 assign mul_22_25_n_1711 = (mul_22_25_n_1718 ^ (mul_22_25_n_1719 ^ mul_22_25_n_1720));
 assign mul_22_25_n_1689 = ((mul_22_25_n_1716 & mul_22_25_n_1717) | (mul_22_25_n_1715 & (mul_22_25_n_1716
    ^ mul_22_25_n_1717)));
 assign mul_22_25_n_1709 = (mul_22_25_n_1715 ^ (mul_22_25_n_1716 ^ mul_22_25_n_1717));
 assign mul_22_25_n_1687 = ((mul_22_25_n_1713 & mul_22_25_n_1714) | (mul_22_25_n_1712 & (mul_22_25_n_1713
    ^ mul_22_25_n_1714)));
 assign mul_22_25_n_1707 = (mul_22_25_n_1712 ^ (mul_22_25_n_1713 ^ mul_22_25_n_1714));
 assign mul_22_25_n_1685 = ((mul_22_25_n_1710 & mul_22_25_n_1711) | (mul_22_25_n_1709 & (mul_22_25_n_1710
    ^ mul_22_25_n_1711)));
 assign mul_22_25_n_1705 = (mul_22_25_n_1709 ^ (mul_22_25_n_1710 ^ mul_22_25_n_1711));
 assign mul_22_25_n_1682 = ((n_148 & n_173) | (n_105 & (n_148 ^ n_173)));
 assign mul_22_25_n_1704 = (n_105 ^ (n_148 ^ n_173));
 assign mul_22_25_n_2293 = ((mul_22_25_n_1704 & n_174) | (mul_22_25_n_1703 & (mul_22_25_n_1704 ^ n_174)));
 assign mul_22_25_n_2253 = (mul_22_25_n_1703 ^ (mul_22_25_n_1704 ^ n_174));
 assign mul_22_25_n_1680 = ((mul_22_25_n_904 & mul_22_25_n_868) | (mul_22_25_n_720 & (mul_22_25_n_904
    ^ mul_22_25_n_868)));
 assign mul_22_25_n_1697 = (mul_22_25_n_720 ^ (mul_22_25_n_904 ^ mul_22_25_n_868));
 assign mul_22_25_n_1679 = ((mul_22_25_n_984 & mul_22_25_n_971) | (mul_22_25_n_805 & (mul_22_25_n_984
    ^ mul_22_25_n_971)));
 assign mul_22_25_n_1696 = (mul_22_25_n_805 ^ (mul_22_25_n_984 ^ mul_22_25_n_971));
 assign mul_22_25_n_1681 = ((mul_22_25_n_1026 & mul_22_25_n_1080) | (mul_22_25_n_1044 & (mul_22_25_n_1026
    ^ mul_22_25_n_1080)));
 assign mul_22_25_n_1698 = (mul_22_25_n_1044 ^ (mul_22_25_n_1026 ^ mul_22_25_n_1080));
 assign mul_22_25_n_1674 = ((mul_22_25_n_782 & mul_22_25_n_872) | (mul_22_25_n_911 & (mul_22_25_n_782
    ^ mul_22_25_n_872)));
 assign mul_22_25_n_1695 = (mul_22_25_n_911 ^ (mul_22_25_n_782 ^ mul_22_25_n_872));
 assign mul_22_25_n_1673 = ((mul_22_25_n_1701 & mul_22_25_n_1702) | (mul_22_25_n_1700 & (mul_22_25_n_1701
    ^ mul_22_25_n_1702)));
 assign mul_22_25_n_1692 = (mul_22_25_n_1700 ^ (mul_22_25_n_1701 ^ mul_22_25_n_1702));
 assign mul_22_25_n_1672 = ((mul_22_25_n_1698 & mul_22_25_n_1699) | (mul_22_25_n_1697 & (mul_22_25_n_1698
    ^ mul_22_25_n_1699)));
 assign mul_22_25_n_1690 = (mul_22_25_n_1697 ^ (mul_22_25_n_1698 ^ mul_22_25_n_1699));
 assign mul_22_25_n_1668 = ((mul_22_25_n_1695 & mul_22_25_n_1696) | (mul_22_25_n_1694 & (mul_22_25_n_1695
    ^ mul_22_25_n_1696)));
 assign mul_22_25_n_1688 = (mul_22_25_n_1694 ^ (mul_22_25_n_1695 ^ mul_22_25_n_1696));
 assign mul_22_25_n_1667 = ((mul_22_25_n_1692 & mul_22_25_n_1693) | (mul_22_25_n_1691 & (mul_22_25_n_1692
    ^ mul_22_25_n_1693)));
 assign mul_22_25_n_1686 = (mul_22_25_n_1691 ^ (mul_22_25_n_1692 ^ mul_22_25_n_1693));
 assign mul_22_25_n_1665 = ((mul_22_25_n_1689 & mul_22_25_n_1690) | (mul_22_25_n_1688 & (mul_22_25_n_1689
    ^ mul_22_25_n_1690)));
 assign mul_22_25_n_1684 = (mul_22_25_n_1688 ^ (mul_22_25_n_1689 ^ mul_22_25_n_1690));
 assign mul_22_25_n_1662 = ((n_58 & n_149) | (n_175 & (n_58 ^ n_149)));
 assign mul_22_25_n_1683 = (n_175 ^ (n_58 ^ n_149));
 assign mul_22_25_n_2294 = ((mul_22_25_n_1683 & n_59) | (mul_22_25_n_1682 & (mul_22_25_n_1683 ^ n_59)));
 assign mul_22_25_n_2254 = (mul_22_25_n_1682 ^ (mul_22_25_n_1683 ^ n_59));
 assign mul_22_25_n_1659 = ((mul_22_25_n_795 & mul_22_25_n_1087) | (mul_22_25_n_1101 & (mul_22_25_n_795
    ^ mul_22_25_n_1087)));
 assign mul_22_25_n_1676 = (mul_22_25_n_1101 ^ (mul_22_25_n_795 ^ mul_22_25_n_1087));
 assign mul_22_25_n_1658 = ((mul_22_25_n_901 & mul_22_25_n_703) | (mul_22_25_n_919 & (mul_22_25_n_901
    ^ mul_22_25_n_703)));
 assign mul_22_25_n_1675 = (mul_22_25_n_919 ^ (mul_22_25_n_901 ^ mul_22_25_n_703));
 assign mul_22_25_n_1661 = ((mul_22_25_n_926 & mul_22_25_n_701) | (mul_22_25_n_927 & (mul_22_25_n_926
    ^ mul_22_25_n_701)));
 assign mul_22_25_n_1678 = (mul_22_25_n_927 ^ (mul_22_25_n_926 ^ mul_22_25_n_701));
 assign mul_22_25_n_1660 = ((mul_22_25_n_793 & mul_22_25_n_935) | (mul_22_25_n_699 & (mul_22_25_n_793
    ^ mul_22_25_n_935)));
 assign mul_22_25_n_1677 = (mul_22_25_n_699 ^ (mul_22_25_n_793 ^ mul_22_25_n_935));
 assign mul_22_25_n_1654 = ((mul_22_25_n_1681 & mul_22_25_n_910) | (mul_22_25_n_1680 & (mul_22_25_n_1681
    ^ mul_22_25_n_910)));
 assign mul_22_25_n_1671 = (mul_22_25_n_1680 ^ (mul_22_25_n_1681 ^ mul_22_25_n_910));
 assign mul_22_25_n_1651 = ((mul_22_25_n_1678 & mul_22_25_n_1679) | (mul_22_25_n_1677 & (mul_22_25_n_1678
    ^ mul_22_25_n_1679)));
 assign mul_22_25_n_1670 = (mul_22_25_n_1677 ^ (mul_22_25_n_1678 ^ mul_22_25_n_1679));
 assign mul_22_25_n_1650 = ((mul_22_25_n_1675 & mul_22_25_n_1676) | (mul_22_25_n_1674 & (mul_22_25_n_1675
    ^ mul_22_25_n_1676)));
 assign mul_22_25_n_1669 = (mul_22_25_n_1674 ^ (mul_22_25_n_1675 ^ mul_22_25_n_1676));
 assign mul_22_25_n_1647 = ((mul_22_25_n_1672 & mul_22_25_n_1673) | (mul_22_25_n_1671 & (mul_22_25_n_1672
    ^ mul_22_25_n_1673)));
 assign mul_22_25_n_1666 = (mul_22_25_n_1671 ^ (mul_22_25_n_1672 ^ mul_22_25_n_1673));
 assign mul_22_25_n_1646 = ((mul_22_25_n_1669 & mul_22_25_n_1670) | (mul_22_25_n_1668 & (mul_22_25_n_1669
    ^ mul_22_25_n_1670)));
 assign mul_22_25_n_1664 = (mul_22_25_n_1668 ^ (mul_22_25_n_1669 ^ mul_22_25_n_1670));
 assign mul_22_25_n_1643 = ((mul_22_25_n_1666 & mul_22_25_n_1667) | (mul_22_25_n_1665 & (mul_22_25_n_1666
    ^ mul_22_25_n_1667)));
 assign mul_22_25_n_1663 = (mul_22_25_n_1665 ^ (mul_22_25_n_1666 ^ mul_22_25_n_1667));
 assign mul_22_25_n_2295 = ((n_133 & n_109) | (mul_22_25_n_1662 & (n_133 ^ n_109)));
 assign mul_22_25_n_2255 = (mul_22_25_n_1662 ^ (n_133 ^ n_109));
 assign mul_22_25_n_1641 = ((mul_22_25_n_745 & mul_22_25_n_707) | (mul_22_25_n_693 & (mul_22_25_n_745
    ^ mul_22_25_n_707)));
 assign mul_22_25_n_1655 = (mul_22_25_n_693 ^ (mul_22_25_n_745 ^ mul_22_25_n_707));
 assign mul_22_25_n_1640 = ((mul_22_25_n_691 & mul_22_25_n_790) | (mul_22_25_n_798 & (mul_22_25_n_691
    ^ mul_22_25_n_790)));
 assign mul_22_25_n_1656 = (mul_22_25_n_798 ^ (mul_22_25_n_691 ^ mul_22_25_n_790));
 assign mul_22_25_n_1642 = ((mul_22_25_n_828 & mul_22_25_n_1091) | (mul_22_25_n_862 & (mul_22_25_n_828
    ^ mul_22_25_n_1091)));
 assign mul_22_25_n_1657 = (mul_22_25_n_862 ^ (mul_22_25_n_828 ^ mul_22_25_n_1091));
 assign mul_22_25_n_1634 = ((mul_22_25_n_1134 & mul_22_25_n_689) | (mul_22_25_n_1661 & (mul_22_25_n_1134
    ^ mul_22_25_n_689)));
 assign mul_22_25_n_1653 = (mul_22_25_n_1661 ^ (mul_22_25_n_1134 ^ mul_22_25_n_689));
 assign mul_22_25_n_1635 = ((mul_22_25_n_1659 & mul_22_25_n_1660) | (mul_22_25_n_1658 & (mul_22_25_n_1659
    ^ mul_22_25_n_1660)));
 assign mul_22_25_n_1652 = (mul_22_25_n_1658 ^ (mul_22_25_n_1659 ^ mul_22_25_n_1660));
 assign mul_22_25_n_1632 = ((mul_22_25_n_1656 & mul_22_25_n_1657) | (mul_22_25_n_1655 & (mul_22_25_n_1656
    ^ mul_22_25_n_1657)));
 assign mul_22_25_n_1649 = (mul_22_25_n_1655 ^ (mul_22_25_n_1656 ^ mul_22_25_n_1657));
 assign mul_22_25_n_1629 = ((mul_22_25_n_1653 & mul_22_25_n_1654) | (mul_22_25_n_1652 & (mul_22_25_n_1653
    ^ mul_22_25_n_1654)));
 assign mul_22_25_n_1648 = (mul_22_25_n_1652 ^ (mul_22_25_n_1653 ^ mul_22_25_n_1654));
 assign mul_22_25_n_1627 = ((mul_22_25_n_1650 & mul_22_25_n_1651) | (mul_22_25_n_1649 & (mul_22_25_n_1650
    ^ mul_22_25_n_1651)));
 assign mul_22_25_n_1645 = (mul_22_25_n_1649 ^ (mul_22_25_n_1650 ^ mul_22_25_n_1651));
 assign mul_22_25_n_1625 = ((mul_22_25_n_1647 & mul_22_25_n_1648) | (mul_22_25_n_1646 & (mul_22_25_n_1647
    ^ mul_22_25_n_1648)));
 assign mul_22_25_n_1644 = (mul_22_25_n_1646 ^ (mul_22_25_n_1647 ^ mul_22_25_n_1648));
 assign mul_22_25_n_2296 = ((n_131 & n_107) | (n_134 & (n_131 ^ n_107)));
 assign mul_22_25_n_2256 = (n_134 ^ (n_131 ^ n_107));
 assign mul_22_25_n_1624 = ((mul_22_25_n_1037 & mul_22_25_n_1094) | (mul_22_25_n_1043 & (mul_22_25_n_1037
    ^ mul_22_25_n_1094)));
 assign mul_22_25_n_1637 = (mul_22_25_n_1043 ^ (mul_22_25_n_1037 ^ mul_22_25_n_1094));
 assign mul_22_25_n_1623 = ((mul_22_25_n_1052 & mul_22_25_n_717) | (mul_22_25_n_751 & (mul_22_25_n_1052
    ^ mul_22_25_n_717)));
 assign mul_22_25_n_1639 = (mul_22_25_n_751 ^ (mul_22_25_n_1052 ^ mul_22_25_n_717));
 assign mul_22_25_n_1622 = ((mul_22_25_n_972 & mul_22_25_n_1065) | (mul_22_25_n_1049 & (mul_22_25_n_972
    ^ mul_22_25_n_1065)));
 assign mul_22_25_n_1638 = (mul_22_25_n_1049 ^ (mul_22_25_n_972 ^ mul_22_25_n_1065));
 assign mul_22_25_n_1618 = ((mul_22_25_n_1046 & mul_22_25_n_954) | (mul_22_25_n_1135 & (mul_22_25_n_1046
    ^ mul_22_25_n_954)));
 assign mul_22_25_n_1636 = (mul_22_25_n_1135 ^ (mul_22_25_n_1046 ^ mul_22_25_n_954));
 assign mul_22_25_n_1617 = ((mul_22_25_n_1641 & mul_22_25_n_1642) | (mul_22_25_n_1640 & (mul_22_25_n_1641
    ^ mul_22_25_n_1642)));
 assign mul_22_25_n_1633 = (mul_22_25_n_1640 ^ (mul_22_25_n_1641 ^ mul_22_25_n_1642));
 assign mul_22_25_n_1616 = ((mul_22_25_n_1638 & mul_22_25_n_1639) | (mul_22_25_n_1637 & (mul_22_25_n_1638
    ^ mul_22_25_n_1639)));
 assign mul_22_25_n_1631 = (mul_22_25_n_1637 ^ (mul_22_25_n_1638 ^ mul_22_25_n_1639));
 assign mul_22_25_n_1612 = ((mul_22_25_n_1635 & mul_22_25_n_1636) | (mul_22_25_n_1634 & (mul_22_25_n_1635
    ^ mul_22_25_n_1636)));
 assign mul_22_25_n_1630 = (mul_22_25_n_1634 ^ (mul_22_25_n_1635 ^ mul_22_25_n_1636));
 assign mul_22_25_n_1611 = ((mul_22_25_n_1632 & mul_22_25_n_1633) | (mul_22_25_n_1631 & (mul_22_25_n_1632
    ^ mul_22_25_n_1633)));
 assign mul_22_25_n_1628 = (mul_22_25_n_1631 ^ (mul_22_25_n_1632 ^ mul_22_25_n_1633));
 assign mul_22_25_n_1608 = ((mul_22_25_n_1629 & mul_22_25_n_1630) | (mul_22_25_n_1628 & (mul_22_25_n_1629
    ^ mul_22_25_n_1630)));
 assign mul_22_25_n_1626 = (mul_22_25_n_1628 ^ (mul_22_25_n_1629 ^ mul_22_25_n_1630));
 assign mul_22_25_n_2297 = ((n_51 & n_108) | (n_132 & (n_51 ^ n_108)));
 assign mul_22_25_n_2257 = (n_132 ^ (n_51 ^ n_108));
 assign mul_22_25_n_1607 = ((mul_22_25_n_711 & mul_22_25_n_1041) | (mul_22_25_n_1038 & (mul_22_25_n_711
    ^ mul_22_25_n_1041)));
 assign mul_22_25_n_1621 = (mul_22_25_n_1038 ^ (mul_22_25_n_711 ^ mul_22_25_n_1041));
 assign mul_22_25_n_1606 = ((mul_22_25_n_1036 & mul_22_25_n_823) | (mul_22_25_n_898 & (mul_22_25_n_1036
    ^ mul_22_25_n_823)));
 assign mul_22_25_n_1620 = (mul_22_25_n_898 ^ (mul_22_25_n_1036 ^ mul_22_25_n_823));
 assign mul_22_25_n_1605 = ((mul_22_25_n_1014 & mul_22_25_n_1033) | (mul_22_25_n_1031 & (mul_22_25_n_1014
    ^ mul_22_25_n_1033)));
 assign mul_22_25_n_1619 = (mul_22_25_n_1031 ^ (mul_22_25_n_1014 ^ mul_22_25_n_1033));
 assign mul_22_25_n_1600 = ((mul_22_25_n_1624 & mul_22_25_n_1) | (mul_22_25_n_1623 & (mul_22_25_n_1624
    ^ mul_22_25_n_1)));
 assign mul_22_25_n_1615 = (mul_22_25_n_1623 ^ (mul_22_25_n_1624 ^ mul_22_25_n_1));
 assign mul_22_25_n_1599 = ((mul_22_25_n_1621 & mul_22_25_n_1622) | (mul_22_25_n_1620 & (mul_22_25_n_1621
    ^ mul_22_25_n_1622)));
 assign mul_22_25_n_1614 = (mul_22_25_n_1620 ^ (mul_22_25_n_1621 ^ mul_22_25_n_1622));
 assign mul_22_25_n_1596 = ((mul_22_25_n_1618 & mul_22_25_n_1619) | (mul_22_25_n_1617 & (mul_22_25_n_1618
    ^ mul_22_25_n_1619)));
 assign mul_22_25_n_1613 = (mul_22_25_n_1617 ^ (mul_22_25_n_1618 ^ mul_22_25_n_1619));
 assign mul_22_25_n_1595 = ((mul_22_25_n_1615 & mul_22_25_n_1616) | (mul_22_25_n_1614 & (mul_22_25_n_1615
    ^ mul_22_25_n_1616)));
 assign mul_22_25_n_1610 = (mul_22_25_n_1614 ^ (mul_22_25_n_1615 ^ mul_22_25_n_1616));
 assign mul_22_25_n_1592 = ((mul_22_25_n_1612 & mul_22_25_n_1613) | (mul_22_25_n_1611 & (mul_22_25_n_1612
    ^ mul_22_25_n_1613)));
 assign mul_22_25_n_1609 = (mul_22_25_n_1611 ^ (mul_22_25_n_1612 ^ mul_22_25_n_1613));
 assign mul_22_25_n_2298 = ((n_78 & n_156) | (n_52 & (n_78 ^ n_156)));
 assign mul_22_25_n_2258 = (n_52 ^ (n_78 ^ n_156));
 assign mul_22_25_n_1591 = ((mul_22_25_n_763 & mul_22_25_n_1090) | (mul_22_25_n_1088 & (mul_22_25_n_763
    ^ mul_22_25_n_1090)));
 assign mul_22_25_n_1603 = (mul_22_25_n_1088 ^ (mul_22_25_n_763 ^ mul_22_25_n_1090));
 assign mul_22_25_n_1590 = ((mul_22_25_n_952 & mul_22_25_n_1021) | (mul_22_25_n_949 & (mul_22_25_n_952
    ^ mul_22_25_n_1021)));
 assign mul_22_25_n_1602 = (mul_22_25_n_949 ^ (mul_22_25_n_952 ^ mul_22_25_n_1021));
 assign mul_22_25_n_1589 = ((mul_22_25_n_1025 & mul_22_25_n_1002) | (mul_22_25_n_831 & (mul_22_25_n_1025
    ^ mul_22_25_n_1002)));
 assign mul_22_25_n_1604 = (mul_22_25_n_831 ^ (mul_22_25_n_1025 ^ mul_22_25_n_1002));
 assign mul_22_25_n_1585 = ((mul_22_25_n_1136 & mul_22_25_n_1018) | (mul_22_25_n_1607 & (mul_22_25_n_1136
    ^ mul_22_25_n_1018)));
 assign mul_22_25_n_1601 = (mul_22_25_n_1607 ^ (mul_22_25_n_1136 ^ mul_22_25_n_1018));
 assign mul_22_25_n_1584 = ((mul_22_25_n_1605 & mul_22_25_n_1606) | (mul_22_25_n_1604 & (mul_22_25_n_1605
    ^ mul_22_25_n_1606)));
 assign mul_22_25_n_1598 = (mul_22_25_n_1604 ^ (mul_22_25_n_1605 ^ mul_22_25_n_1606));
 assign mul_22_25_n_1581 = ((mul_22_25_n_1602 & mul_22_25_n_1603) | (mul_22_25_n_1601 & (mul_22_25_n_1602
    ^ mul_22_25_n_1603)));
 assign mul_22_25_n_1597 = (mul_22_25_n_1601 ^ (mul_22_25_n_1602 ^ mul_22_25_n_1603));
 assign mul_22_25_n_1580 = ((mul_22_25_n_1599 & mul_22_25_n_1600) | (mul_22_25_n_1598 & (mul_22_25_n_1599
    ^ mul_22_25_n_1600)));
 assign mul_22_25_n_1594 = (mul_22_25_n_1598 ^ (mul_22_25_n_1599 ^ mul_22_25_n_1600));
 assign mul_22_25_n_1577 = ((mul_22_25_n_1596 & mul_22_25_n_1597) | (mul_22_25_n_1595 & (mul_22_25_n_1596
    ^ mul_22_25_n_1597)));
 assign mul_22_25_n_1593 = (mul_22_25_n_1595 ^ (mul_22_25_n_1596 ^ mul_22_25_n_1597));
 assign mul_22_25_n_2299 = ((n_154 & n_116) | (n_79 & (n_154 ^ n_116)));
 assign mul_22_25_n_2259 = (n_79 ^ (n_154 ^ n_116));
 assign mul_22_25_n_1576 = ((mul_22_25_n_1099 & mul_22_25_n_1010) | (mul_22_25_n_957 & (mul_22_25_n_1099
    ^ mul_22_25_n_1010)));
 assign mul_22_25_n_1588 = (mul_22_25_n_957 ^ (mul_22_25_n_1099 ^ mul_22_25_n_1010));
 assign mul_22_25_n_1575 = ((mul_22_25_n_1001 & mul_22_25_n_873) | (mul_22_25_n_1007 & (mul_22_25_n_1001
    ^ mul_22_25_n_873)));
 assign mul_22_25_n_1587 = (mul_22_25_n_1007 ^ (mul_22_25_n_1001 ^ mul_22_25_n_873));
 assign mul_22_25_n_1571 = ((mul_22_25_n_830 & mul_22_25_n_1006) | (mul_22_25_n_1138 & (mul_22_25_n_830
    ^ mul_22_25_n_1006)));
 assign mul_22_25_n_1586 = (mul_22_25_n_1138 ^ (mul_22_25_n_830 ^ mul_22_25_n_1006));
 assign mul_22_25_n_1570 = ((mul_22_25_n_1590 & mul_22_25_n_1591) | (mul_22_25_n_1589 & (mul_22_25_n_1590
    ^ mul_22_25_n_1591)));
 assign mul_22_25_n_1583 = (mul_22_25_n_1589 ^ (mul_22_25_n_1590 ^ mul_22_25_n_1591));
 assign mul_22_25_n_1567 = ((mul_22_25_n_1587 & mul_22_25_n_1588) | (mul_22_25_n_1586 & (mul_22_25_n_1587
    ^ mul_22_25_n_1588)));
 assign mul_22_25_n_1582 = (mul_22_25_n_1586 ^ (mul_22_25_n_1587 ^ mul_22_25_n_1588));
 assign mul_22_25_n_1566 = ((mul_22_25_n_1584 & mul_22_25_n_1585) | (mul_22_25_n_1583 & (mul_22_25_n_1584
    ^ mul_22_25_n_1585)));
 assign mul_22_25_n_1579 = (mul_22_25_n_1583 ^ (mul_22_25_n_1584 ^ mul_22_25_n_1585));
 assign mul_22_25_n_1563 = ((mul_22_25_n_1581 & mul_22_25_n_1582) | (mul_22_25_n_1580 & (mul_22_25_n_1581
    ^ mul_22_25_n_1582)));
 assign mul_22_25_n_1578 = (mul_22_25_n_1580 ^ (mul_22_25_n_1581 ^ mul_22_25_n_1582));
 assign mul_22_25_n_2300 = ((n_114 & n_113) | (n_155 & (n_114 ^ n_113)));
 assign mul_22_25_n_2260 = (n_155 ^ (n_114 ^ n_113));
 assign mul_22_25_n_1562 = ((mul_22_25_n_1024 & mul_22_25_n_1081) | (mul_22_25_n_1000 & (mul_22_25_n_1024
    ^ mul_22_25_n_1081)));
 assign mul_22_25_n_1574 = (mul_22_25_n_1000 ^ (mul_22_25_n_1024 ^ mul_22_25_n_1081));
 assign mul_22_25_n_1561 = ((mul_22_25_n_744 & mul_22_25_n_814) | (mul_22_25_n_804 & (mul_22_25_n_744
    ^ mul_22_25_n_814)));
 assign mul_22_25_n_1572 = (mul_22_25_n_804 ^ (mul_22_25_n_744 ^ mul_22_25_n_814));
 assign mul_22_25_n_1560 = ((mul_22_25_n_964 & mul_22_25_n_996) | (mul_22_25_n_754 & (mul_22_25_n_964
    ^ mul_22_25_n_996)));
 assign mul_22_25_n_1573 = (mul_22_25_n_754 ^ (mul_22_25_n_964 ^ mul_22_25_n_996));
 assign mul_22_25_n_1556 = ((mul_22_25_n_1576 & mul_22_25_n_1137) | (mul_22_25_n_1575 & (mul_22_25_n_1576
    ^ mul_22_25_n_1137)));
 assign mul_22_25_n_1569 = (mul_22_25_n_1575 ^ (mul_22_25_n_1576 ^ mul_22_25_n_1137));
 assign mul_22_25_n_1554 = ((mul_22_25_n_1573 & mul_22_25_n_1574) | (mul_22_25_n_1572 & (mul_22_25_n_1573
    ^ mul_22_25_n_1574)));
 assign mul_22_25_n_1568 = (mul_22_25_n_1572 ^ (mul_22_25_n_1573 ^ mul_22_25_n_1574));
 assign mul_22_25_n_1552 = ((mul_22_25_n_1570 & mul_22_25_n_1571) | (mul_22_25_n_1569 & (mul_22_25_n_1570
    ^ mul_22_25_n_1571)));
 assign mul_22_25_n_1565 = (mul_22_25_n_1569 ^ (mul_22_25_n_1570 ^ mul_22_25_n_1571));
 assign mul_22_25_n_1550 = ((mul_22_25_n_1567 & mul_22_25_n_1568) | (mul_22_25_n_1566 & (mul_22_25_n_1567
    ^ mul_22_25_n_1568)));
 assign mul_22_25_n_1564 = (mul_22_25_n_1566 ^ (mul_22_25_n_1567 ^ mul_22_25_n_1568));
 assign mul_22_25_n_2301 = ((n_142 & n_111) | (n_115 & (n_142 ^ n_111)));
 assign mul_22_25_n_2261 = (n_115 ^ (n_142 ^ n_111));
 assign mul_22_25_n_1548 = ((mul_22_25_n_1042 & mul_22_25_n_860) | (mul_22_25_n_1035 & (mul_22_25_n_1042
    ^ mul_22_25_n_860)));
 assign mul_22_25_n_1558 = (mul_22_25_n_1035 ^ (mul_22_25_n_1042 ^ mul_22_25_n_860));
 assign mul_22_25_n_1549 = ((mul_22_25_n_985 & mul_22_25_n_990) | (mul_22_25_n_921 & (mul_22_25_n_985
    ^ mul_22_25_n_990)));
 assign mul_22_25_n_1559 = (mul_22_25_n_921 ^ (mul_22_25_n_985 ^ mul_22_25_n_990));
 assign mul_22_25_n_1544 = ((mul_22_25_n_0 & mul_22_25_n_951) | (mul_22_25_n_1562 & (mul_22_25_n_0 ^
    mul_22_25_n_951)));
 assign mul_22_25_n_1557 = (mul_22_25_n_1562 ^ (mul_22_25_n_0 ^ mul_22_25_n_951));
 assign mul_22_25_n_1542 = ((mul_22_25_n_1560 & mul_22_25_n_1561) | (mul_22_25_n_1559 & (mul_22_25_n_1560
    ^ mul_22_25_n_1561)));
 assign mul_22_25_n_1555 = (mul_22_25_n_1559 ^ (mul_22_25_n_1560 ^ mul_22_25_n_1561));
 assign mul_22_25_n_1541 = ((mul_22_25_n_1557 & mul_22_25_n_1558) | (mul_22_25_n_1556 & (mul_22_25_n_1557
    ^ mul_22_25_n_1558)));
 assign mul_22_25_n_1553 = (mul_22_25_n_1556 ^ (mul_22_25_n_1557 ^ mul_22_25_n_1558));
 assign mul_22_25_n_1538 = ((mul_22_25_n_1554 & mul_22_25_n_1555) | (mul_22_25_n_1553 & (mul_22_25_n_1554
    ^ mul_22_25_n_1555)));
 assign mul_22_25_n_1551 = (mul_22_25_n_1553 ^ (mul_22_25_n_1554 ^ mul_22_25_n_1555));
 assign mul_22_25_n_2302 = ((n_45 & n_112) | (n_143 & (n_45 ^ n_112)));
 assign mul_22_25_n_2262 = (n_143 ^ (n_45 ^ n_112));
 assign mul_22_25_n_1537 = ((mul_22_25_n_826 & mul_22_25_n_1089) | (mul_22_25_n_708 & (mul_22_25_n_826
    ^ mul_22_25_n_1089)));
 assign mul_22_25_n_1547 = (mul_22_25_n_708 ^ (mul_22_25_n_826 ^ mul_22_25_n_1089));
 assign mul_22_25_n_1536 = ((mul_22_25_n_1030 & mul_22_25_n_979) | (mul_22_25_n_884 & (mul_22_25_n_1030
    ^ mul_22_25_n_979)));
 assign mul_22_25_n_1546 = (mul_22_25_n_884 ^ (mul_22_25_n_1030 ^ mul_22_25_n_979));
 assign mul_22_25_n_1533 = ((mul_22_25_n_975 & mul_22_25_n_977) | (mul_22_25_n_1141 & (mul_22_25_n_975
    ^ mul_22_25_n_977)));
 assign mul_22_25_n_1545 = (mul_22_25_n_1141 ^ (mul_22_25_n_975 ^ mul_22_25_n_977));
 assign mul_22_25_n_1531 = ((mul_22_25_n_1548 & mul_22_25_n_1549) | (mul_22_25_n_1547 & (mul_22_25_n_1548
    ^ mul_22_25_n_1549)));
 assign mul_22_25_n_1543 = (mul_22_25_n_1547 ^ (mul_22_25_n_1548 ^ mul_22_25_n_1549));
 assign mul_22_25_n_1529 = ((mul_22_25_n_1545 & mul_22_25_n_1546) | (mul_22_25_n_1544 & (mul_22_25_n_1545
    ^ mul_22_25_n_1546)));
 assign mul_22_25_n_1540 = (mul_22_25_n_1544 ^ (mul_22_25_n_1545 ^ mul_22_25_n_1546));
 assign mul_22_25_n_1527 = ((mul_22_25_n_1542 & mul_22_25_n_1543) | (mul_22_25_n_1541 & (mul_22_25_n_1542
    ^ mul_22_25_n_1543)));
 assign mul_22_25_n_1539 = (mul_22_25_n_1541 ^ (mul_22_25_n_1542 ^ mul_22_25_n_1543));
 assign mul_22_25_n_2264 = ((n_50 & n_101) | (n_46 & (n_50 ^ n_101)));
 assign mul_22_25_n_2263 = (n_46 ^ (n_50 ^ n_101));
 assign asc001_26_ = (mul_22_25_n_1336 ^ mul_22_25_n_1416);
 assign asc001_47_ = (mul_22_25_n_1325 ^ mul_22_25_n_1511);
 assign asc001_49_ = ~(mul_22_25_n_10 ^ mul_22_25_n_1500);
 assign mul_22_25_n_1511 = ~(mul_22_25_n_1311 | (mul_22_25_n_1506 & mul_22_25_n_1300));
 assign asc001_46_ = ~(mul_22_25_n_1323 ^ mul_22_25_n_1506);
 assign asc001_45_ = ~(mul_22_25_n_1327 ^ mul_22_25_n_1505);
 assign asc001_43_ = ~(mul_22_25_n_1421 ^ mul_22_25_n_1504);
 assign asc001_39_ = ~(mul_22_25_n_1418 ^ mul_22_25_n_1498);
 assign mul_22_25_n_1506 = ~(mul_22_25_n_1347 & (mul_22_25_n_1494 | mul_22_25_n_1345));
 assign mul_22_25_n_1505 = ~(mul_22_25_n_1310 & (mul_22_25_n_1494 | mul_22_25_n_1315));
 assign mul_22_25_n_1504 = ~(mul_22_25_n_1386 & (mul_22_25_n_1493 | mul_22_25_n_1384));
 assign asc001_44_ = (mul_22_25_n_1326 ^ mul_22_25_n_1494);
 assign asc001_42_ = (mul_22_25_n_1420 ^ mul_22_25_n_1493);
 assign asc001_41_ = ~(mul_22_25_n_1422 ^ mul_22_25_n_1492);
 assign mul_22_25_n_1500 = ~(mul_22_25_n_1320 | (mul_22_25_n_1491 & mul_22_25_n_1309));
 assign asc001_48_ = ~(mul_22_25_n_1334 ^ mul_22_25_n_1491);
 assign mul_22_25_n_1498 = ~(mul_22_25_n_1396 & (mul_22_25_n_1489 | mul_22_25_n_1390));
 assign asc001_38_ = ~(mul_22_25_n_1417 ^ mul_22_25_n_1489);
 assign asc001_37_ = ~(mul_22_25_n_1408 ^ mul_22_25_n_1488);
 assign asc001_35_ = ~(mul_22_25_n_1461 ^ mul_22_25_n_1487);
 assign mul_22_25_n_1494 = ~(mul_22_25_n_1455 | (mul_22_25_n_1483 & mul_22_25_n_1433));
 assign mul_22_25_n_1493 = ~(mul_22_25_n_1430 | (mul_22_25_n_1483 & mul_22_25_n_1426));
 assign mul_22_25_n_1492 = (~mul_22_25_n_1383 | (mul_22_25_n_1483 & mul_22_25_n_1394));
 assign mul_22_25_n_1491 = ~(mul_22_25_n_1471 & (mul_22_25_n_1477 & (mul_22_25_n_1482 | mul_22_25_n_1451)));
 assign asc001_40_ = ~(mul_22_25_n_1419 ^ mul_22_25_n_1483);
 assign mul_22_25_n_1489 = ~(mul_22_25_n_1432 | (mul_22_25_n_1481 & mul_22_25_n_1427));
 assign mul_22_25_n_1488 = (~mul_22_25_n_1389 | (mul_22_25_n_1481 & mul_22_25_n_12));
 assign mul_22_25_n_1487 = ~(mul_22_25_n_1448 & (mul_22_25_n_1480 | mul_22_25_n_1450));
 assign asc001_36_ = ~(mul_22_25_n_1406 ^ mul_22_25_n_1481);
 assign asc001_34_ = ~(mul_22_25_n_1460 ^ mul_22_25_n_1480);
 assign asc001_33_ = ~(mul_22_25_n_1459 ^ mul_22_25_n_1479);
 assign mul_22_25_n_1483 = ~(mul_22_25_n_1482 & (mul_22_25_n_1475 | mul_22_25_n_1472));
 assign mul_22_25_n_1482 = ~(mul_22_25_n_1447 | (mul_22_25_n_1431 | (mul_22_25_n_1476 & mul_22_25_n_1435)));
 assign mul_22_25_n_1481 = ~(~mul_22_25_n_1476 & (mul_22_25_n_1475 | mul_22_25_n_1469));
 assign mul_22_25_n_1480 = (~mul_22_25_n_1468 & (mul_22_25_n_1475 | mul_22_25_n_1457));
 assign mul_22_25_n_1479 = ~(mul_22_25_n_1444 & (mul_22_25_n_1475 | mul_22_25_n_1445));
 assign asc001_32_ = ~(mul_22_25_n_1458 ^ mul_22_25_n_1475);
 assign mul_22_25_n_1477 = (mul_22_25_n_1451 | (mul_22_25_n_1472 | mul_22_25_n_1475));
 assign mul_22_25_n_1476 = ~(mul_22_25_n_1452 & (mul_22_25_n_1473 & (mul_22_25_n_1449 | mul_22_25_n_1448)));
 assign mul_22_25_n_1475 = ~(mul_22_25_n_1470 | (mul_22_25_n_1364 & mul_22_25_n_1454));
 assign asc001_31_ = ~(mul_22_25_n_1405 ^ mul_22_25_n_1467);
 assign mul_22_25_n_1473 = ~(mul_22_25_n_1468 & mul_22_25_n_1462);
 assign mul_22_25_n_1472 = ~(~mul_22_25_n_1469 & mul_22_25_n_1435);
 assign mul_22_25_n_1471 = ~(mul_22_25_n_1360 | (mul_22_25_n_1350 | (mul_22_25_n_1455 & mul_22_25_n_1354)));
 assign mul_22_25_n_1470 = ~(mul_22_25_n_1456 & (mul_22_25_n_1463 & (mul_22_25_n_1381 | mul_22_25_n_1436)));
 assign mul_22_25_n_1469 = ~(~mul_22_25_n_1457 & mul_22_25_n_1462);
 assign mul_22_25_n_1468 = ~(mul_22_25_n_1453 & (mul_22_25_n_1442 | mul_22_25_n_1444));
 assign mul_22_25_n_1467 = ~(mul_22_25_n_1401 | (mul_22_25_n_1443 & mul_22_25_n_1400));
 assign asc001_27_ = ~(mul_22_25_n_1367 ^ mul_22_25_n_1438);
 assign asc001_30_ = ~(mul_22_25_n_1411 ^ mul_22_25_n_1443);
 assign asc001_29_ = ~(mul_22_25_n_1410 ^ mul_22_25_n_1437);
 assign mul_22_25_n_1463 = ~(mul_22_25_n_1369 & mul_22_25_n_1454);
 assign mul_22_25_n_1462 = ~(mul_22_25_n_1449 | mul_22_25_n_1450);
 assign mul_22_25_n_1461 = ~(mul_22_25_n_1452 & ~mul_22_25_n_1449);
 assign mul_22_25_n_1460 = ~(mul_22_25_n_1450 | ~mul_22_25_n_1448);
 assign mul_22_25_n_1459 = ~(~mul_22_25_n_1442 & mul_22_25_n_1453);
 assign mul_22_25_n_1458 = ~(~mul_22_25_n_1444 | mul_22_25_n_1445);
 assign mul_22_25_n_1457 = (mul_22_25_n_1442 | mul_22_25_n_1445);
 assign mul_22_25_n_1456 = ~(mul_22_25_n_1423 | (mul_22_25_n_1403 | (mul_22_25_n_1434 & mul_22_25_n_1424)));
 assign mul_22_25_n_1455 = ~(mul_22_25_n_1392 & (mul_22_25_n_1446 & (mul_22_25_n_1385 | mul_22_25_n_1386)));
 assign mul_22_25_n_1447 = (mul_22_25_n_1432 & mul_22_25_n_1428);
 assign mul_22_25_n_1446 = ~(mul_22_25_n_1430 & mul_22_25_n_1425);
 assign mul_22_25_n_1454 = ~(mul_22_25_n_1436 | mul_22_25_n_1371);
 assign mul_22_25_n_1453 = ~(mul_22_25_n_2248 & mul_22_25_n_2287);
 assign mul_22_25_n_1452 = ~(mul_22_25_n_2250 & mul_22_25_n_2289);
 assign mul_22_25_n_1451 = ~(mul_22_25_n_1354 & mul_22_25_n_1433);
 assign mul_22_25_n_1450 = ~(mul_22_25_n_2249 | mul_22_25_n_2288);
 assign mul_22_25_n_1449 = ~(mul_22_25_n_2250 | mul_22_25_n_2289);
 assign mul_22_25_n_1448 = ~(mul_22_25_n_2249 & mul_22_25_n_2288);
 assign asc001_23_ = ~(mul_22_25_n_1339 ^ mul_22_25_n_1407);
 assign asc001_25_ = ~(mul_22_25_n_1341 ^ mul_22_25_n_13);
 assign asc001_28_ = ~(mul_22_25_n_1409 ^ mul_22_25_n_1415);
 assign mul_22_25_n_1438 = ~(mul_22_25_n_1318 | (mul_22_25_n_1416 & mul_22_25_n_1317));
 assign mul_22_25_n_1437 = ~(mul_22_25_n_1397 | (mul_22_25_n_1414 & mul_22_25_n_1395));
 assign mul_22_25_n_1445 = ~(mul_22_25_n_2247 | mul_22_25_n_2286);
 assign mul_22_25_n_1444 = ~(mul_22_25_n_2247 & mul_22_25_n_2286);
 assign mul_22_25_n_1443 = ~(~mul_22_25_n_1434 & (mul_22_25_n_1415 | mul_22_25_n_1429));
 assign mul_22_25_n_1442 = ~(mul_22_25_n_2248 | mul_22_25_n_2287);
 assign mul_22_25_n_1431 = ~(mul_22_25_n_1402 & (mul_22_25_n_1387 | mul_22_25_n_1396));
 assign mul_22_25_n_1436 = ~(mul_22_25_n_1424 & ~mul_22_25_n_1429);
 assign mul_22_25_n_1435 = (mul_22_25_n_1428 & mul_22_25_n_1427);
 assign mul_22_25_n_1434 = (~mul_22_25_n_1404 | (mul_22_25_n_15 & mul_22_25_n_1397));
 assign mul_22_25_n_1433 = (mul_22_25_n_1425 & mul_22_25_n_1426);
 assign mul_22_25_n_1432 = ~(mul_22_25_n_1393 & (mul_22_25_n_1388 | mul_22_25_n_1389));
 assign mul_22_25_n_1430 = ~(mul_22_25_n_1391 & (mul_22_25_n_1399 | mul_22_25_n_1383));
 assign mul_22_25_n_1423 = (mul_22_25_n_1398 & mul_22_25_n_1401);
 assign mul_22_25_n_1422 = ~(~mul_22_25_n_1399 & mul_22_25_n_1391);
 assign mul_22_25_n_1429 = ~(mul_22_25_n_15 & mul_22_25_n_1395);
 assign mul_22_25_n_1428 = ~(mul_22_25_n_1387 | mul_22_25_n_1390);
 assign mul_22_25_n_1427 = ~(mul_22_25_n_1388 | ~mul_22_25_n_12);
 assign mul_22_25_n_1421 = ~(~mul_22_25_n_1385 & mul_22_25_n_1392);
 assign mul_22_25_n_1420 = ~(mul_22_25_n_1386 & ~mul_22_25_n_1384);
 assign mul_22_25_n_1426 = ~(mul_22_25_n_1399 | ~mul_22_25_n_1394);
 assign mul_22_25_n_1425 = ~(mul_22_25_n_1385 | mul_22_25_n_1384);
 assign mul_22_25_n_1419 = ~(mul_22_25_n_1394 & mul_22_25_n_1383);
 assign mul_22_25_n_1418 = ~(mul_22_25_n_1402 & ~mul_22_25_n_1387);
 assign mul_22_25_n_1417 = ~(mul_22_25_n_1390 | ~mul_22_25_n_1396);
 assign mul_22_25_n_1424 = (mul_22_25_n_1398 & mul_22_25_n_1400);
 assign mul_22_25_n_1415 = ~mul_22_25_n_1414;
 assign asc001_21_ = ~(mul_22_25_n_1337 ^ mul_22_25_n_11);
 assign asc001_24_ = ~(mul_22_25_n_1340 ^ mul_22_25_n_1375);
 assign mul_22_25_n_1411 = ~(~mul_22_25_n_1401 & mul_22_25_n_1400);
 assign mul_22_25_n_1410 = (mul_22_25_n_15 & mul_22_25_n_1404);
 assign mul_22_25_n_1409 = ~(mul_22_25_n_1397 | ~mul_22_25_n_1395);
 assign mul_22_25_n_1408 = ~(mul_22_25_n_1393 & ~mul_22_25_n_1388);
 assign mul_22_25_n_1407 = ~(mul_22_25_n_1298 & (mul_22_25_n_1376 | mul_22_25_n_1303));
 assign mul_22_25_n_1406 = ~(mul_22_25_n_12 & mul_22_25_n_1389);
 assign mul_22_25_n_1405 = ~(mul_22_25_n_1403 | ~mul_22_25_n_1398);
 assign mul_22_25_n_1416 = ~(mul_22_25_n_1353 & (mul_22_25_n_1375 | mul_22_25_n_1344));
 assign mul_22_25_n_1414 = ~(mul_22_25_n_1381 & (mul_22_25_n_1375 | mul_22_25_n_1371));
 assign mul_22_25_n_1404 = ~(mul_22_25_n_2244 & mul_22_25_n_2283);
 assign mul_22_25_n_1403 = ~(mul_22_25_n_1379 | mul_22_25_n_1380);
 assign mul_22_25_n_1402 = ~(mul_22_25_n_2254 & mul_22_25_n_2293);
 assign mul_22_25_n_1401 = ~(mul_22_25_n_1377 | mul_22_25_n_1378);
 assign mul_22_25_n_1400 = ~(mul_22_25_n_1377 & mul_22_25_n_1378);
 assign mul_22_25_n_1399 = ~(mul_22_25_n_2256 | mul_22_25_n_2295);
 assign mul_22_25_n_1398 = ~(mul_22_25_n_1379 & mul_22_25_n_1380);
 assign mul_22_25_n_1397 = ~(mul_22_25_n_1382 | mul_22_25_n_1346);
 assign mul_22_25_n_1396 = ~(mul_22_25_n_2253 & mul_22_25_n_2292);
 assign mul_22_25_n_1395 = ~(mul_22_25_n_1382 & mul_22_25_n_1346);
 assign mul_22_25_n_1394 = ~(mul_22_25_n_1372 & mul_22_25_n_1373);
 assign mul_22_25_n_1393 = ~(mul_22_25_n_2252 & mul_22_25_n_2291);
 assign mul_22_25_n_1392 = ~(mul_22_25_n_2258 & mul_22_25_n_2297);
 assign mul_22_25_n_1391 = ~(mul_22_25_n_2256 & mul_22_25_n_2295);
 assign mul_22_25_n_1390 = ~(mul_22_25_n_2253 | mul_22_25_n_2292);
 assign mul_22_25_n_1389 = ~(mul_22_25_n_2251 & mul_22_25_n_2290);
 assign mul_22_25_n_1388 = ~(mul_22_25_n_2252 | mul_22_25_n_2291);
 assign mul_22_25_n_1387 = ~(mul_22_25_n_2254 | mul_22_25_n_2293);
 assign mul_22_25_n_1386 = ~(mul_22_25_n_2257 & mul_22_25_n_2296);
 assign mul_22_25_n_1385 = ~(mul_22_25_n_2258 | mul_22_25_n_2297);
 assign mul_22_25_n_1384 = ~(mul_22_25_n_2257 | mul_22_25_n_2296);
 assign mul_22_25_n_1383 = (mul_22_25_n_1372 | mul_22_25_n_1373);
 assign mul_22_25_n_1382 = ~mul_22_25_n_2243;
 assign mul_22_25_n_1380 = ~mul_22_25_n_2285;
 assign mul_22_25_n_1379 = ~mul_22_25_n_2246;
 assign mul_22_25_n_1378 = ~mul_22_25_n_2284;
 assign mul_22_25_n_1377 = ~mul_22_25_n_2245;
 assign asc001_20_ = ~(mul_22_25_n_1342 ^ mul_22_25_n_1366);
 assign mul_22_25_n_1381 = ~(mul_22_25_n_1363 | (mul_22_25_n_1370 | (mul_22_25_n_1362 & mul_22_25_n_1318)));
 assign mul_22_25_n_1376 = ~(mul_22_25_n_1351 | (mul_22_25_n_1366 & mul_22_25_n_1333));
 assign mul_22_25_n_1375 = ~(mul_22_25_n_1364 | mul_22_25_n_1369);
 assign mul_22_25_n_1373 = ~mul_22_25_n_2294;
 assign mul_22_25_n_1372 = ~mul_22_25_n_2255;
 assign mul_22_25_n_1370 = ~(mul_22_25_n_1353 | mul_22_25_n_1365);
 assign mul_22_25_n_1371 = (mul_22_25_n_1365 | mul_22_25_n_1344);
 assign asc001_19_ = ~(mul_22_25_n_1335 ^ mul_22_25_n_1359);
 assign mul_22_25_n_1369 = ~(mul_22_25_n_1361 & (mul_22_25_n_1349 & (mul_22_25_n_1358 | mul_22_25_n_1352)));
 assign mul_22_25_n_1367 = ~(mul_22_25_n_1363 | ~mul_22_25_n_1362);
 assign mul_22_25_n_1366 = ~(mul_22_25_n_1357 & mul_22_25_n_1358);
 assign mul_22_25_n_1365 = ~(mul_22_25_n_1362 & mul_22_25_n_1317);
 assign mul_22_25_n_1364 = ~(mul_22_25_n_1357 | mul_22_25_n_1352);
 assign mul_22_25_n_1363 = ~(mul_22_25_n_1348 | mul_22_25_n_1295);
 assign mul_22_25_n_1362 = ~(mul_22_25_n_1348 & mul_22_25_n_1295);
 assign mul_22_25_n_1361 = ~(mul_22_25_n_1351 & mul_22_25_n_1343);
 assign mul_22_25_n_1360 = ~(mul_22_25_n_1347 | mul_22_25_n_1331);
 assign mul_22_25_n_1359 = ~(mul_22_25_n_1275 & (mul_22_25_n_1330 | mul_22_25_n_1274));
 assign mul_22_25_n_1358 = ~(mul_22_25_n_1329 | (mul_22_25_n_1308 | (mul_22_25_n_1269 & mul_22_25_n_1332)));
 assign mul_22_25_n_1357 = ~(mul_22_25_n_1332 & (mul_22_25_n_1263 & mul_22_25_n_1286));
 assign asc001_18_ = ~(mul_22_25_n_1278 ^ mul_22_25_n_1330);
 assign asc001_17_ = ~(mul_22_25_n_1265 ^ mul_22_25_n_1324);
 assign mul_22_25_n_1350 = (~mul_22_25_n_1321 | (mul_22_25_n_1304 & mul_22_25_n_1311));
 assign mul_22_25_n_1349 = (~mul_22_25_n_1319 & (mul_22_25_n_1297 | mul_22_25_n_1298));
 assign mul_22_25_n_1354 = ~(mul_22_25_n_1331 | mul_22_25_n_1345);
 assign mul_22_25_n_1353 = ~(mul_22_25_n_1322 | (mul_22_25_n_1313 & mul_22_25_n_1314));
 assign mul_22_25_n_1352 = ~(mul_22_25_n_1343 & mul_22_25_n_1333);
 assign mul_22_25_n_1351 = ~(mul_22_25_n_1307 & (mul_22_25_n_1299 | mul_22_25_n_1302));
 assign mul_22_25_n_1348 = ~mul_22_25_n_2242;
 assign mul_22_25_n_1346 = ~mul_22_25_n_2282;
 assign mul_22_25_n_1347 = (~mul_22_25_n_1306 & (mul_22_25_n_1316 | mul_22_25_n_1310));
 assign mul_22_25_n_1342 = ~(~mul_22_25_n_1305 & mul_22_25_n_1302);
 assign mul_22_25_n_1341 = ~(mul_22_25_n_1322 | ~mul_22_25_n_1313);
 assign mul_22_25_n_1340 = ~(mul_22_25_n_1314 | ~mul_22_25_n_1312);
 assign mul_22_25_n_1339 = (mul_22_25_n_1297 | mul_22_25_n_1319);
 assign mul_22_25_n_1338 = ~(~mul_22_25_n_1303 & mul_22_25_n_1298);
 assign mul_22_25_n_1337 = ~(mul_22_25_n_1307 & ~mul_22_25_n_1299);
 assign mul_22_25_n_1336 = ~(mul_22_25_n_1318 | ~mul_22_25_n_1317);
 assign mul_22_25_n_1335 = ~(~mul_22_25_n_1308 & mul_22_25_n_1301);
 assign mul_22_25_n_1345 = (mul_22_25_n_1316 | mul_22_25_n_1315);
 assign mul_22_25_n_1344 = ~(mul_22_25_n_1313 & mul_22_25_n_1312);
 assign mul_22_25_n_1343 = ~(mul_22_25_n_1297 | mul_22_25_n_1303);
 assign mul_22_25_n_1334 = ~(~mul_22_25_n_1320 & mul_22_25_n_1309);
 assign mul_22_25_n_1329 = ~(~mul_22_25_n_1301 | mul_22_25_n_1275);
 assign asc001_16_ = ~(mul_22_25_n_1266 ^ mul_22_25_n_1286);
 assign mul_22_25_n_1327 = (mul_22_25_n_1316 | mul_22_25_n_1306);
 assign mul_22_25_n_1333 = ~(mul_22_25_n_1299 | mul_22_25_n_1305);
 assign mul_22_25_n_1326 = ~(mul_22_25_n_1310 & ~mul_22_25_n_1315);
 assign mul_22_25_n_1332 = ~(~mul_22_25_n_1301 | mul_22_25_n_1274);
 assign mul_22_25_n_1325 = ~(mul_22_25_n_1304 & mul_22_25_n_1321);
 assign mul_22_25_n_1331 = ~(mul_22_25_n_1304 & mul_22_25_n_1300);
 assign mul_22_25_n_1324 = (~mul_22_25_n_1256 | (mul_22_25_n_1286 & mul_22_25_n_9));
 assign mul_22_25_n_1323 = ~(~mul_22_25_n_1311 & mul_22_25_n_1300);
 assign mul_22_25_n_1330 = ~(mul_22_25_n_1269 | (mul_22_25_n_1286 & mul_22_25_n_1263));
 assign mul_22_25_n_1322 = ~(mul_22_25_n_1289 | mul_22_25_n_1290);
 assign mul_22_25_n_1321 = ~(mul_22_25_n_2262 & mul_22_25_n_2301);
 assign mul_22_25_n_1320 = ~(mul_22_25_n_1294 | mul_22_25_n_1292);
 assign mul_22_25_n_1319 = ~(mul_22_25_n_1285 | mul_22_25_n_1281);
 assign mul_22_25_n_1318 = ~(mul_22_25_n_1293 | mul_22_25_n_1291);
 assign mul_22_25_n_1317 = ~(mul_22_25_n_1293 & mul_22_25_n_1291);
 assign mul_22_25_n_1316 = ~(mul_22_25_n_2260 | mul_22_25_n_2299);
 assign mul_22_25_n_1315 = ~(mul_22_25_n_2259 | mul_22_25_n_2298);
 assign mul_22_25_n_1314 = ~(mul_22_25_n_1287 | mul_22_25_n_1288);
 assign mul_22_25_n_1313 = ~(mul_22_25_n_1289 & mul_22_25_n_1290);
 assign mul_22_25_n_1312 = ~(mul_22_25_n_1287 & mul_22_25_n_1288);
 assign mul_22_25_n_1311 = ~(mul_22_25_n_1282 | mul_22_25_n_1283);
 assign mul_22_25_n_1310 = ~(mul_22_25_n_2259 & mul_22_25_n_2298);
 assign asc001_15_ = ~(mul_22_25_n_1264 ^ mul_22_25_n_1280);
 assign mul_22_25_n_1309 = ~(mul_22_25_n_1294 & mul_22_25_n_1292);
 assign mul_22_25_n_1308 = ~(mul_22_25_n_1284 | n_93);
 assign mul_22_25_n_1307 = ~(mul_22_25_n_2236 & mul_22_25_n_2275);
 assign mul_22_25_n_1306 = (mul_22_25_n_2260 & mul_22_25_n_2299);
 assign mul_22_25_n_1305 = ~(mul_22_25_n_2235 | mul_22_25_n_2274);
 assign mul_22_25_n_1304 = (mul_22_25_n_2262 | mul_22_25_n_2301);
 assign mul_22_25_n_1303 = ~(mul_22_25_n_2237 | mul_22_25_n_2276);
 assign mul_22_25_n_1302 = ~(mul_22_25_n_2235 & mul_22_25_n_2274);
 assign mul_22_25_n_1301 = ~(mul_22_25_n_1284 & n_93);
 assign mul_22_25_n_1300 = ~(mul_22_25_n_1282 & mul_22_25_n_1283);
 assign mul_22_25_n_1299 = ~(mul_22_25_n_2236 | mul_22_25_n_2275);
 assign mul_22_25_n_1298 = ~(mul_22_25_n_2237 & mul_22_25_n_2276);
 assign mul_22_25_n_1297 = (mul_22_25_n_1285 & mul_22_25_n_1281);
 assign mul_22_25_n_1295 = ~mul_22_25_n_2281;
 assign mul_22_25_n_1294 = ~mul_22_25_n_2263;
 assign mul_22_25_n_1293 = ~mul_22_25_n_2241;
 assign mul_22_25_n_1292 = ~mul_22_25_n_2302;
 assign mul_22_25_n_1291 = ~mul_22_25_n_2280;
 assign mul_22_25_n_1290 = ~mul_22_25_n_2279;
 assign mul_22_25_n_1289 = ~mul_22_25_n_2240;
 assign mul_22_25_n_1288 = ~mul_22_25_n_2278;
 assign mul_22_25_n_1287 = ~mul_22_25_n_2239;
 assign mul_22_25_n_1286 = ~(mul_22_25_n_1276 & (mul_22_25_n_1277 & (mul_22_25_n_1234 | mul_22_25_n_1271)));
 assign mul_22_25_n_1285 = ~mul_22_25_n_2238;
 assign mul_22_25_n_1284 = ~mul_22_25_n_2234;
 assign mul_22_25_n_1283 = ~mul_22_25_n_2300;
 assign mul_22_25_n_1282 = ~mul_22_25_n_2261;
 assign mul_22_25_n_1281 = ~mul_22_25_n_2277;
 assign mul_22_25_n_1280 = ~(n_47 | (mul_22_25_n_1273 & n_84));
 assign asc001_14_ = ~(mul_22_25_n_1259 ^ mul_22_25_n_1273);
 assign mul_22_25_n_1278 = ~(~mul_22_25_n_1275 | mul_22_25_n_1274);
 assign mul_22_25_n_1277 = ~(mul_22_25_n_1261 | (n_81 | (mul_22_25_n_1270 & mul_22_25_n_1262)));
 assign mul_22_25_n_1276 = (mul_22_25_n_1239 | mul_22_25_n_1271);
 assign mul_22_25_n_1275 = ~(n_94 & n_86);
 assign mul_22_25_n_1274 = ~(n_94 | n_86);
 assign mul_22_25_n_1273 = ~(~mul_22_25_n_1270 & (mul_22_25_n_1242 | mul_22_25_n_1267));
 assign asc001_13_ = ~(mul_22_25_n_1260 ^ mul_22_25_n_1247);
 assign mul_22_25_n_1271 = ~(~mul_22_25_n_1267 & mul_22_25_n_1262);
 assign mul_22_25_n_1270 = ~(n_55 & (n_54 | n_88));
 assign mul_22_25_n_1269 = ~(n_95 & (n_57 | mul_22_25_n_1256));
 assign mul_22_25_n_1268 = ~mul_22_25_n_2273;
 assign mul_22_25_n_1266 = ~(mul_22_25_n_9 & mul_22_25_n_1256);
 assign mul_22_25_n_1265 = ~(~n_57 & n_95);
 assign mul_22_25_n_1267 = (n_54 | n_85);
 assign mul_22_25_n_1264 = ~(n_83 | n_81);
 assign mul_22_25_n_1261 = ~(n_83 | ~n_47);
 assign mul_22_25_n_1260 = ~(n_54 | ~n_55);
 assign mul_22_25_n_1259 = ~(n_84 & ~n_47);
 assign mul_22_25_n_1263 = ~(n_57 | ~mul_22_25_n_9);
 assign mul_22_25_n_1262 = ~(~n_84 | n_83);
 assign mul_22_25_n_1258 = ~(mul_22_25_n_2232 & mul_22_25_n_2271);
 assign mul_22_25_n_1257 = ~(mul_22_25_n_1245 | mul_22_25_n_1246);
 assign mul_22_25_n_1256 = ~(n_96 & n_135);
 assign mul_22_25_n_1255 = ~(mul_22_25_n_2232 | mul_22_25_n_2271);
 assign mul_22_25_n_1254 = ~(mul_22_25_n_2228 | mul_22_25_n_2267);
 assign asc001_11_ = (mul_22_25_n_1229 ^ mul_22_25_n_1241);
 assign asc001_12_ = ~(mul_22_25_n_1240 ^ mul_22_25_n_1242);
 assign mul_22_25_n_1247 = (n_88 & (mul_22_25_n_1242 | n_85));
 assign mul_22_25_n_1253 = ~(mul_22_25_n_2228 & mul_22_25_n_2267);
 assign mul_22_25_n_1252 = ~(mul_22_25_n_1243 & mul_22_25_n_1244);
 assign mul_22_25_n_1251 = ~(mul_22_25_n_1243 | mul_22_25_n_1244);
 assign mul_22_25_n_1250 = (mul_22_25_n_1245 & mul_22_25_n_1246);
 assign mul_22_25_n_1246 = ~mul_22_25_n_2269;
 assign mul_22_25_n_1245 = ~mul_22_25_n_2230;
 assign mul_22_25_n_1244 = ~mul_22_25_n_2268;
 assign mul_22_25_n_1243 = ~mul_22_25_n_2229;
 assign mul_22_25_n_1242 = (mul_22_25_n_1234 & mul_22_25_n_1239);
 assign mul_22_25_n_1241 = ~(n_89 & (mul_22_25_n_1236 | n_56));
 assign mul_22_25_n_1240 = ~(~n_88 | n_85);
 assign mul_22_25_n_1239 = ~(mul_22_25_n_1230 | (n_90 | (n_91 & mul_22_25_n_1231)));
 assign mul_22_25_n_1238 = ~(mul_22_25_n_1514 & mul_22_25_n_1516);
 assign mul_22_25_n_1237 = ~(mul_22_25_n_1514 | mul_22_25_n_1516);
 assign mul_22_25_n_1236 = ~(n_123 | n_91);
 assign asc001_9_ = ~(n_65 ^ n_122);
 assign mul_22_25_n_1234 = ~(n_123 & mul_22_25_n_1231);
 assign mul_22_25_n_1233 = ~(mul_22_25_n_1222 & (mul_22_25_n_1221 | mul_22_25_n_1212));
 assign mul_22_25_n_1230 = ~(n_87 | n_89);
 assign mul_22_25_n_1232 = ~(mul_22_25_n_1216 | mul_22_25_n_1221);
 assign mul_22_25_n_1231 = ~(n_87 | n_56);
 assign mul_22_25_n_1229 = ~(n_87 | n_90);
 assign mul_22_25_n_1228 = ~(n_56 | ~n_89);
 assign mul_22_25_n_1227 = ~(mul_22_25_n_1221 | ~mul_22_25_n_1222);
 assign mul_22_25_n_1226 = ~(mul_22_25_n_1219 | mul_22_25_n_1220);
 assign mul_22_25_n_1225 = ~(mul_22_25_n_2227 & mul_22_25_n_1518);
 assign mul_22_25_n_1224 = (mul_22_25_n_1219 & mul_22_25_n_1220);
 assign mul_22_25_n_1223 = ~(mul_22_25_n_2227 | mul_22_25_n_1518);
 assign mul_22_25_n_1222 = ~(mul_22_25_n_2226 & mul_22_25_n_2266);
 assign mul_22_25_n_1221 = ~(mul_22_25_n_2226 | mul_22_25_n_2266);
 assign mul_22_25_n_1220 = ~mul_22_25_n_1517;
 assign mul_22_25_n_1219 = ~mul_22_25_n_1515;
 assign asc001_8_ = ~(mul_22_25_n_1215 ^ mul_22_25_n_1214);
 assign mul_22_25_n_1217 = (mul_22_25_n_1216 & mul_22_25_n_1212);
 assign mul_22_25_n_1216 = ~(~mul_22_25_n_1214 & mul_22_25_n_1211);
 assign mul_22_25_n_1215 = (mul_22_25_n_1211 & mul_22_25_n_1212);
 assign mul_22_25_n_1214 = ~(mul_22_25_n_1209 | (mul_22_25_n_1208 | (mul_22_25_n_1197 & mul_22_25_n_1206)));
 assign asc001_7_ = (mul_22_25_n_1205 ^ mul_22_25_n_1207);
 assign mul_22_25_n_1212 = ~(mul_22_25_n_1519 & mul_22_25_n_1521);
 assign mul_22_25_n_1211 = (mul_22_25_n_1519 | mul_22_25_n_1521);
 assign asc001_6_ = ~(mul_22_25_n_1199 ^ mul_22_25_n_1204);
 assign mul_22_25_n_1209 = ~(mul_22_25_n_1203 & (mul_22_25_n_1201 | mul_22_25_n_1202));
 assign mul_22_25_n_1208 = (mul_22_25_n_1196 & mul_22_25_n_1206);
 assign mul_22_25_n_1207 = ~(mul_22_25_n_1202 & (mul_22_25_n_1199 | mul_22_25_n_1200));
 assign mul_22_25_n_1206 = ~(mul_22_25_n_1201 | mul_22_25_n_1200);
 assign mul_22_25_n_1205 = ~(~mul_22_25_n_1203 | mul_22_25_n_1201);
 assign mul_22_25_n_1204 = ~(mul_22_25_n_1200 | ~mul_22_25_n_1202);
 assign mul_22_25_n_1203 = ~(mul_22_25_n_1520 & mul_22_25_n_1523);
 assign mul_22_25_n_1202 = ~(mul_22_25_n_1522 & mul_22_25_n_2265);
 assign mul_22_25_n_1201 = ~(mul_22_25_n_1520 | mul_22_25_n_1523);
 assign mul_22_25_n_1200 = ~(mul_22_25_n_1522 | mul_22_25_n_2265);
 assign asc001_5_ = ~(mul_22_25_n_1191 ^ mul_22_25_n_1195);
 assign mul_22_25_n_1199 = ~(mul_22_25_n_1196 | mul_22_25_n_1197);
 assign mul_22_25_n_1197 = ~(mul_22_25_n_1194 & (mul_22_25_n_1188 | mul_22_25_n_1193));
 assign mul_22_25_n_1196 = ~(mul_22_25_n_1189 | mul_22_25_n_1193);
 assign mul_22_25_n_1195 = ~(mul_22_25_n_1193 | ~mul_22_25_n_1194);
 assign mul_22_25_n_1194 = ~(mul_22_25_n_1524 & mul_22_25_n_1526);
 assign mul_22_25_n_1193 = ~(mul_22_25_n_1524 | mul_22_25_n_1526);
 assign asc001_4_ = ~(mul_22_25_n_1186 ^ mul_22_25_n_1190);
 assign mul_22_25_n_1191 = (mul_22_25_n_1189 & mul_22_25_n_1188);
 assign mul_22_25_n_1190 = ~(mul_22_25_n_1188 & mul_22_25_n_1187);
 assign mul_22_25_n_1189 = ~(mul_22_25_n_1186 & mul_22_25_n_1187);
 assign mul_22_25_n_1188 = ~(mul_22_25_n_1161 & mul_22_25_n_1525);
 assign mul_22_25_n_1187 = (mul_22_25_n_1161 | mul_22_25_n_1525);
 assign asc001_3_ = (mul_22_25_n_1182 ^ mul_22_25_n_1183);
 assign mul_22_25_n_1186 = ~(mul_22_25_n_1184 & (mul_22_25_n_1180 & (mul_22_25_n_1181 | mul_22_25_n_1178)));
 assign mul_22_25_n_1184 = ~(mul_22_25_n_1133 & ~mul_22_25_n_1181);
 assign mul_22_25_n_1183 = ~(~mul_22_25_n_1180 | mul_22_25_n_1181);
 assign mul_22_25_n_1182 = ~(~mul_22_25_n_1133 & mul_22_25_n_1178);
 assign mul_22_25_n_1181 = ~(mul_22_25_n_1169 | mul_22_25_n_1142);
 assign mul_22_25_n_1180 = ~(mul_22_25_n_1169 & mul_22_25_n_1142);
 assign asc001_2_ = ~(mul_22_25_n_1113 ^ mul_22_25_n_1153);
 assign mul_22_25_n_1178 = ~(mul_22_25_n_1143 & mul_22_25_n_1113);
 assign mul_22_25_n_1177 = ~(mul_22_25_n_1116 ^ mul_22_25_n_686);
 assign mul_22_25_n_1176 = (mul_22_25_n_1118 ^ mul_22_25_n_909);
 assign mul_22_25_n_1175 = ~(mul_22_25_n_1120 ^ mul_22_25_n_908);
 assign mul_22_25_n_1174 = ~(mul_22_25_n_1124 ^ mul_22_25_n_1131);
 assign mul_22_25_n_1173 = ~(mul_22_25_n_1152 & (mul_22_25_n_914 | mul_22_25_n_688));
 assign mul_22_25_n_1172 = ~(mul_22_25_n_1121 ^ mul_22_25_n_1114);
 assign mul_22_25_n_1171 = (mul_22_25_n_1128 ^ mul_22_25_n_1115);
 assign mul_22_25_n_1170 = (mul_22_25_n_1119 ^ mul_22_25_n_1132);
 assign mul_22_25_n_1168 = (mul_22_25_n_1130 ^ mul_22_25_n_659);
 assign mul_22_25_n_1167 = (mul_22_25_n_1123 ^ mul_22_25_n_685);
 assign mul_22_25_n_1166 = (mul_22_25_n_1126 ^ mul_22_25_n_661);
 assign mul_22_25_n_1165 = (mul_22_25_n_658 ^ mul_22_25_n_1117);
 assign mul_22_25_n_1164 = (mul_22_25_n_663 ^ mul_22_25_n_1129);
 assign mul_22_25_n_1163 = (mul_22_25_n_1125 ^ mul_22_25_n_657);
 assign mul_22_25_n_1162 = (mul_22_25_n_662 ^ mul_22_25_n_1127);
 assign mul_22_25_n_1169 = (mul_22_25_n_660 ^ mul_22_25_n_1122);
 assign mul_22_25_n_1160 = ~(mul_22_25_n_658 | mul_22_25_n_1117);
 assign mul_22_25_n_1159 = ~(mul_22_25_n_657 | mul_22_25_n_1125);
 assign mul_22_25_n_1158 = ~(mul_22_25_n_685 | mul_22_25_n_1123);
 assign mul_22_25_n_1157 = ~(mul_22_25_n_661 | mul_22_25_n_1126);
 assign mul_22_25_n_1156 = ~(mul_22_25_n_662 | mul_22_25_n_1127);
 assign mul_22_25_n_1155 = ~(mul_22_25_n_659 | mul_22_25_n_1130);
 assign mul_22_25_n_1154 = ~(mul_22_25_n_663 | mul_22_25_n_1129);
 assign mul_22_25_n_1161 = ~(mul_22_25_n_660 | mul_22_25_n_1122);
 assign mul_22_25_n_1153 = ~(mul_22_25_n_1143 & ~mul_22_25_n_1133);
 assign asc001_1_ = ~(mul_22_25_n_1113 | (mul_22_25_n_687 & mul_22_25_n_508));
 assign mul_22_25_n_1150 = ~(mul_22_25_n_909 | mul_22_25_n_1118);
 assign mul_22_25_n_1149 = ~(mul_22_25_n_1132 | mul_22_25_n_1119);
 assign mul_22_25_n_1148 = ~(mul_22_25_n_1120 | ~mul_22_25_n_908);
 assign mul_22_25_n_1147 = ~(mul_22_25_n_1121 | ~mul_22_25_n_1114);
 assign mul_22_25_n_1146 = ~(mul_22_25_n_1115 | mul_22_25_n_1128);
 assign mul_22_25_n_1145 = ~(mul_22_25_n_1124 | ~mul_22_25_n_1131);
 assign mul_22_25_n_1144 = ~(mul_22_25_n_1116 | ~mul_22_25_n_686);
 assign mul_22_25_n_1152 = ~(mul_22_25_n_914 & mul_22_25_n_688);
 assign mul_22_25_n_1141 = ~mul_22_25_n_0;
 assign mul_22_25_n_1140 = ~mul_22_25_n_1139;
 assign mul_22_25_n_1138 = ~mul_22_25_n_1137;
 assign mul_22_25_n_1136 = ~mul_22_25_n_1;
 assign mul_22_25_n_1135 = ~mul_22_25_n_1134;
 assign mul_22_25_n_1112 = ~((mul_22_25_n_362 | mul_22_25_n_134) & (mul_22_25_n_617 | mul_22_25_n_124));
 assign mul_22_25_n_1111 = ~((mul_22_25_n_349 | mul_22_25_n_263) & (mul_22_25_n_602 | mul_22_25_n_374));
 assign mul_22_25_n_1110 = ~((mul_22_25_n_351 | mul_22_25_n_545) & (mul_22_25_n_596 | mul_22_25_n_542));
 assign mul_22_25_n_1109 = ~((mul_22_25_n_353 | mul_22_25_n_395) & (mul_22_25_n_610 | mul_22_25_n_399));
 assign mul_22_25_n_1108 = ~((mul_22_25_n_356 | mul_22_25_n_554) & (mul_22_25_n_600 | mul_22_25_n_515));
 assign mul_22_25_n_1107 = ~((mul_22_25_n_356 | mul_22_25_n_386) & (mul_22_25_n_600 | mul_22_25_n_302));
 assign mul_22_25_n_1106 = ~((mul_22_25_n_358 | mul_22_25_n_220) & (mul_22_25_n_613 | mul_22_25_n_219));
 assign mul_22_25_n_1105 = ~((mul_22_25_n_350 | mul_22_25_n_285) & (mul_22_25_n_606 | mul_22_25_n_424));
 assign mul_22_25_n_1104 = ~((mul_22_25_n_359 | mul_22_25_n_202) & (mul_22_25_n_614 | mul_22_25_n_192));
 assign mul_22_25_n_1103 = ~((mul_22_25_n_355 | mul_22_25_n_460) & (mul_22_25_n_598 | mul_22_25_n_372));
 assign mul_22_25_n_1102 = ~((mul_22_25_n_353 | mul_22_25_n_476) & (mul_22_25_n_610 | mul_22_25_n_448));
 assign mul_22_25_n_1101 = ~((mul_22_25_n_350 | mul_22_25_n_518) & (mul_22_25_n_606 | mul_22_25_n_487));
 assign mul_22_25_n_1100 = ~((mul_22_25_n_352 | mul_22_25_n_512) & (mul_22_25_n_604 | mul_22_25_n_521));
 assign mul_22_25_n_1099 = ~((mul_22_25_n_362 | mul_22_25_n_133) & (mul_22_25_n_617 | mul_22_25_n_135));
 assign mul_22_25_n_1098 = ~((mul_22_25_n_358 | mul_22_25_n_215) & (mul_22_25_n_613 | mul_22_25_n_216));
 assign mul_22_25_n_1097 = ~((mul_22_25_n_354 | mul_22_25_n_318) & (mul_22_25_n_612 | mul_22_25_n_270));
 assign mul_22_25_n_1096 = ~((mul_22_25_n_356 | mul_22_25_n_477) & (mul_22_25_n_600 | mul_22_25_n_466));
 assign mul_22_25_n_1095 = ~((mul_22_25_n_353 | mul_22_25_n_579) & (mul_22_25_n_610 | mul_22_25_n_388));
 assign mul_22_25_n_1094 = ~(mul_22_25_n_622 | (mul_22_25_n_607 & mul_22_25_n_565));
 assign mul_22_25_n_1093 = ~((mul_22_25_n_350 | mul_22_25_n_272) & (mul_22_25_n_606 | mul_22_25_n_370));
 assign mul_22_25_n_1092 = ~((mul_22_25_n_352 | mul_22_25_n_384) & (mul_22_25_n_604 | mul_22_25_n_387));
 assign mul_22_25_n_1091 = ~(mul_22_25_n_6 & (mul_22_25_n_608 | mul_22_25_n_569));
 assign mul_22_25_n_1090 = ~(mul_22_25_n_640 | (mul_22_25_n_601 & mul_22_25_n_560));
 assign mul_22_25_n_1089 = ~(mul_22_25_n_2 | (mul_22_25_n_609 & mul_22_25_n_575));
 assign mul_22_25_n_1088 = ~((mul_22_25_n_354 | mul_22_25_n_520) & (mul_22_25_n_612 | mul_22_25_n_494));
 assign mul_22_25_n_1087 = ~(mul_22_25_n_638 | (mul_22_25_n_599 & mul_22_25_n_570));
 assign mul_22_25_n_1086 = ~((mul_22_25_n_355 | mul_22_25_n_496) & (mul_22_25_n_598 | mul_22_25_n_503));
 assign mul_22_25_n_1085 = ~(mul_22_25_n_619 | (mul_22_25_n_595 & mul_22_25_n_559));
 assign mul_22_25_n_1084 = ~(mul_22_25_n_4 & (mul_22_25_n_604 | mul_22_25_n_558));
 assign mul_22_25_n_1083 = ~(mul_22_25_n_620 | (mul_22_25_n_603 & mul_22_25_n_572));
 assign mul_22_25_n_1082 = ~(mul_22_25_n_621 | (mul_22_25_n_597 & mul_22_25_n_566));
 assign mul_22_25_n_1081 = ~(mul_22_25_n_639 | (mul_22_25_n_605 & mul_22_25_n_567));
 assign mul_22_25_n_1080 = ~(mul_22_25_n_5 & (mul_22_25_n_600 | mul_22_25_n_574));
 assign mul_22_25_n_1079 = ~(mul_22_25_n_7 & (mul_22_25_n_598 | mul_22_25_n_564));
 assign mul_22_25_n_1078 = ~((mul_22_25_n_592 & mul_22_25_n_333) | (mul_22_25_n_611 & mul_22_25_n_577));
 assign mul_22_25_n_1077 = ~((mul_22_25_n_358 | mul_22_25_n_332) & (mul_22_25_n_613 | mul_22_25_n_531));
 assign mul_22_25_n_1076 = ~((mul_22_25_n_359 | mul_22_25_n_331) & (mul_22_25_n_614 | mul_22_25_n_507));
 assign mul_22_25_n_1075 = ~((mul_22_25_n_360 | mul_22_25_n_330) & (mul_22_25_n_615 | mul_22_25_n_461));
 assign mul_22_25_n_1074 = ~((mul_22_25_n_361 | mul_22_25_n_329) & (mul_22_25_n_616 | mul_22_25_n_429));
 assign mul_22_25_n_1073 = ~((mul_22_25_n_362 | mul_22_25_n_84) & (mul_22_25_n_617 | mul_22_25_n_161));
 assign mul_22_25_n_1072 = ~((mul_22_25_n_363 | mul_22_25_n_83) & (mul_22_25_n_618 | mul_22_25_n_120));
 assign mul_22_25_n_1071 = ~((mul_22_25_n_363 | mul_22_25_n_108) & (mul_22_25_n_618 | mul_22_25_n_82));
 assign mul_22_25_n_1070 = ~((mul_22_25_n_362 | mul_22_25_n_132) & (mul_22_25_n_617 | mul_22_25_n_81));
 assign mul_22_25_n_1069 = ~((mul_22_25_n_361 | mul_22_25_n_156) & (mul_22_25_n_616 | mul_22_25_n_80));
 assign mul_22_25_n_1068 = ~((mul_22_25_n_357 | mul_22_25_n_281) & (mul_22_25_n_608 | mul_22_25_n_77));
 assign mul_22_25_n_1067 = ~((mul_22_25_n_354 | mul_22_25_n_290) & (mul_22_25_n_612 | mul_22_25_n_75));
 assign mul_22_25_n_1066 = ~((mul_22_25_n_352 | mul_22_25_n_582) & (mul_22_25_n_604 | mul_22_25_n_74));
 assign mul_22_25_n_1065 = ~((mul_22_25_n_362 | mul_22_25_n_122) & (mul_22_25_n_617 | mul_22_25_n_129));
 assign mul_22_25_n_1064 = ~((mul_22_25_n_350 | mul_22_25_n_266) & (mul_22_25_n_606 | mul_22_25_n_73));
 assign mul_22_25_n_1063 = ~((mul_22_25_n_355 | mul_22_25_n_225) & (mul_22_25_n_598 | mul_22_25_n_78));
 assign mul_22_25_n_1062 = ~((mul_22_25_n_356 | mul_22_25_n_371) & (mul_22_25_n_600 | mul_22_25_n_79));
 assign mul_22_25_n_1061 = ~((mul_22_25_n_353 | mul_22_25_n_411) & (mul_22_25_n_610 | mul_22_25_n_85));
 assign mul_22_25_n_1060 = ~((mul_22_25_n_349 | mul_22_25_n_230) & (mul_22_25_n_602 | mul_22_25_n_71));
 assign mul_22_25_n_1059 = ~((mul_22_25_n_360 | mul_22_25_n_173) & (mul_22_25_n_615 | mul_22_25_n_69));
 assign mul_22_25_n_1058 = ~((mul_22_25_n_358 | mul_22_25_n_207) & (mul_22_25_n_613 | mul_22_25_n_68));
 assign mul_22_25_n_1057 = ~((mul_22_25_n_359 | mul_22_25_n_200) & (mul_22_25_n_614 | mul_22_25_n_67));
 assign mul_22_25_n_1056 = ~((mul_22_25_n_349 | mul_22_25_n_473) & (mul_22_25_n_602 | mul_22_25_n_463));
 assign mul_22_25_n_1055 = ~((mul_22_25_n_355 | mul_22_25_n_87) & (mul_22_25_n_598 | mul_22_25_n_300));
 assign mul_22_25_n_1054 = ~((mul_22_25_n_356 | mul_22_25_n_515) & (mul_22_25_n_600 | mul_22_25_n_519));
 assign mul_22_25_n_1053 = ~((mul_22_25_n_353 | mul_22_25_n_412) & (mul_22_25_n_610 | mul_22_25_n_319));
 assign mul_22_25_n_1052 = ~((mul_22_25_n_361 | mul_22_25_n_149) & (mul_22_25_n_616 | mul_22_25_n_146));
 assign mul_22_25_n_1051 = ~((mul_22_25_n_360 | mul_22_25_n_179) & (mul_22_25_n_615 | mul_22_25_n_175));
 assign mul_22_25_n_1050 = ~((mul_22_25_n_353 | mul_22_25_n_399) & (mul_22_25_n_610 | mul_22_25_n_377));
 assign mul_22_25_n_1049 = ~((mul_22_25_n_350 | mul_22_25_n_541) & (mul_22_25_n_606 | mul_22_25_n_523));
 assign mul_22_25_n_1048 = ~((mul_22_25_n_360 | mul_22_25_n_176) & (mul_22_25_n_615 | mul_22_25_n_172));
 assign mul_22_25_n_1047 = ~((mul_22_25_n_358 | mul_22_25_n_213) & (mul_22_25_n_613 | mul_22_25_n_221));
 assign mul_22_25_n_1046 = ~((mul_22_25_n_359 | mul_22_25_n_427) & (mul_22_25_n_614 | mul_22_25_n_184));
 assign mul_22_25_n_1045 = ~((mul_22_25_n_359 | mul_22_25_n_197) & (mul_22_25_n_614 | mul_22_25_n_201));
 assign mul_22_25_n_1044 = ~((mul_22_25_n_363 | mul_22_25_n_110) & (mul_22_25_n_618 | mul_22_25_n_103));
 assign mul_22_25_n_1043 = ~((mul_22_25_n_353 | mul_22_25_n_530) & (mul_22_25_n_610 | mul_22_25_n_491));
 assign mul_22_25_n_1042 = ~((mul_22_25_n_363 | mul_22_25_n_111) & (mul_22_25_n_618 | mul_22_25_n_109));
 assign mul_22_25_n_1041 = ~((mul_22_25_n_354 | mul_22_25_n_494) & (mul_22_25_n_612 | mul_22_25_n_499));
 assign mul_22_25_n_1040 = ~((mul_22_25_n_352 | mul_22_25_n_462) & (mul_22_25_n_604 | mul_22_25_n_469));
 assign mul_22_25_n_1039 = ~((mul_22_25_n_349 | mul_22_25_n_513) & (mul_22_25_n_602 | mul_22_25_n_501));
 assign mul_22_25_n_1038 = ~((mul_22_25_n_362 | mul_22_25_n_139) & (mul_22_25_n_617 | mul_22_25_n_122));
 assign mul_22_25_n_1037 = ~((mul_22_25_n_349 | mul_22_25_n_573) & (mul_22_25_n_602 | mul_22_25_n_551));
 assign mul_22_25_n_1036 = ~((mul_22_25_n_363 | mul_22_25_n_114) & (mul_22_25_n_618 | mul_22_25_n_107));
 assign mul_22_25_n_1035 = ~((mul_22_25_n_359 | mul_22_25_n_483) & (mul_22_25_n_614 | mul_22_25_n_484));
 assign mul_22_25_n_1034 = ~((mul_22_25_n_357 | mul_22_25_n_455) & (mul_22_25_n_608 | mul_22_25_n_443));
 assign mul_22_25_n_1033 = ~((mul_22_25_n_353 | mul_22_25_n_517) & (mul_22_25_n_610 | mul_22_25_n_530));
 assign mul_22_25_n_1032 = ~((mul_22_25_n_349 | mul_22_25_n_393) & (mul_22_25_n_602 | mul_22_25_n_417));
 assign mul_22_25_n_1031 = ~((mul_22_25_n_360 | mul_22_25_n_168) & (mul_22_25_n_615 | mul_22_25_n_165));
 assign mul_22_25_n_1030 = ~((mul_22_25_n_360 | mul_22_25_n_461) & (mul_22_25_n_615 | mul_22_25_n_432));
 assign mul_22_25_n_1029 = ~((mul_22_25_n_357 | mul_22_25_n_506) & (mul_22_25_n_608 | mul_22_25_n_475));
 assign mul_22_25_n_1028 = ~((mul_22_25_n_360 | mul_22_25_n_178) & (mul_22_25_n_615 | mul_22_25_n_167));
 assign mul_22_25_n_1027 = ~((mul_22_25_n_349 | mul_22_25_n_418) & (mul_22_25_n_602 | mul_22_25_n_301));
 assign mul_22_25_n_1026 = ~((mul_22_25_n_349 | mul_22_25_n_529) & (mul_22_25_n_602 | mul_22_25_n_513));
 assign mul_22_25_n_1025 = ~((mul_22_25_n_353 | mul_22_25_n_534) & (mul_22_25_n_610 | mul_22_25_n_517));
 assign mul_22_25_n_1024 = ~((mul_22_25_n_353 | mul_22_25_n_563) & (mul_22_25_n_610 | mul_22_25_n_553));
 assign mul_22_25_n_1023 = ~((mul_22_25_n_359 | mul_22_25_n_201) & (mul_22_25_n_614 | mul_22_25_n_196));
 assign mul_22_25_n_1022 = ~((mul_22_25_n_362 | mul_22_25_n_138) & (mul_22_25_n_617 | mul_22_25_n_131));
 assign mul_22_25_n_1021 = ~((mul_22_25_n_361 | mul_22_25_n_145) & (mul_22_25_n_616 | mul_22_25_n_141));
 assign mul_22_25_n_1020 = ~((mul_22_25_n_351 | mul_22_25_n_181) & (mul_22_25_n_596 | mul_22_25_n_379));
 assign mul_22_25_n_1019 = ~((mul_22_25_n_352 | mul_22_25_n_228) & (mul_22_25_n_604 | mul_22_25_n_288));
 assign mul_22_25_n_1018 = ~((mul_22_25_n_360 | mul_22_25_n_223) & (mul_22_25_n_615 | mul_22_25_n_168));
 assign mul_22_25_n_1017 = ~((mul_22_25_n_352 | mul_22_25_n_414) & (mul_22_25_n_604 | mul_22_25_n_582));
 assign mul_22_25_n_1016 = ~((mul_22_25_n_359 | mul_22_25_n_187) & (mul_22_25_n_614 | mul_22_25_n_190));
 assign mul_22_25_n_1015 = ~((mul_22_25_n_356 | mul_22_25_n_409) & (mul_22_25_n_600 | mul_22_25_n_160));
 assign mul_22_25_n_1014 = ~((mul_22_25_n_359 | mul_22_25_n_426) & (mul_22_25_n_614 | mul_22_25_n_427));
 assign mul_22_25_n_1013 = ~((mul_22_25_n_355 | mul_22_25_n_454) & (mul_22_25_n_598 | mul_22_25_n_436));
 assign mul_22_25_n_1012 = ~((mul_22_25_n_355 | mul_22_25_n_480) & (mul_22_25_n_598 | mul_22_25_n_454));
 assign mul_22_25_n_1011 = ~((mul_22_25_n_352 | mul_22_25_n_398) & (mul_22_25_n_604 | mul_22_25_n_227));
 assign mul_22_25_n_1010 = ~((mul_22_25_n_358 | mul_22_25_n_485) & (mul_22_25_n_613 | mul_22_25_n_486));
 assign mul_22_25_n_1009 = ~((mul_22_25_n_349 | mul_22_25_n_400) & (mul_22_25_n_602 | mul_22_25_n_267));
 assign mul_22_25_n_1008 = ~((mul_22_25_n_354 | mul_22_25_n_270) & (mul_22_25_n_612 | mul_22_25_n_310));
 assign mul_22_25_n_1007 = ~((mul_22_25_n_354 | mul_22_25_n_522) & (mul_22_25_n_612 | mul_22_25_n_520));
 assign mul_22_25_n_1006 = ~((mul_22_25_n_360 | mul_22_25_n_222) & (mul_22_25_n_615 | mul_22_25_n_223));
 assign mul_22_25_n_1005 = ~((mul_22_25_n_351 | mul_22_25_n_498) & (mul_22_25_n_596 | mul_22_25_n_471));
 assign mul_22_25_n_1004 = ~((mul_22_25_n_359 | mul_22_25_n_194) & (mul_22_25_n_614 | mul_22_25_n_197));
 assign mul_22_25_n_1003 = ~((mul_22_25_n_349 | mul_22_25_n_417) & (mul_22_25_n_602 | mul_22_25_n_418));
 assign mul_22_25_n_1002 = ~((mul_22_25_n_363 | mul_22_25_n_117) & (mul_22_25_n_618 | mul_22_25_n_114));
 assign mul_22_25_n_1001 = ~((mul_22_25_n_359 | mul_22_25_n_456) & (mul_22_25_n_614 | mul_22_25_n_457));
 assign mul_22_25_n_1000 = ~((mul_22_25_n_358 | mul_22_25_n_510) & (mul_22_25_n_613 | mul_22_25_n_485));
 assign mul_22_25_n_999 = ~((mul_22_25_n_361 | mul_22_25_n_150) & (mul_22_25_n_616 | mul_22_25_n_151));
 assign mul_22_25_n_998 = ~((mul_22_25_n_354 | mul_22_25_n_115) & (mul_22_25_n_612 | mul_22_25_n_588));
 assign mul_22_25_n_997 = ~((mul_22_25_n_354 | mul_22_25_n_233) & (mul_22_25_n_612 | mul_22_25_n_253));
 assign mul_22_25_n_996 = ~((mul_22_25_n_354 | mul_22_25_n_548) & (mul_22_25_n_612 | mul_22_25_n_522));
 assign mul_22_25_n_995 = ~((mul_22_25_n_361 | mul_22_25_n_151) & (mul_22_25_n_616 | mul_22_25_n_156));
 assign mul_22_25_n_994 = ~((mul_22_25_n_349 | mul_22_25_n_415) & (mul_22_25_n_602 | mul_22_25_n_393));
 assign mul_22_25_n_993 = ~((mul_22_25_n_360 | mul_22_25_n_166) & (mul_22_25_n_615 | mul_22_25_n_173));
 assign mul_22_25_n_992 = ~((mul_22_25_n_358 | mul_22_25_n_221) & (mul_22_25_n_613 | mul_22_25_n_212));
 assign mul_22_25_n_991 = ~((mul_22_25_n_352 | mul_22_25_n_434) & (mul_22_25_n_604 | mul_22_25_n_435));
 assign mul_22_25_n_990 = ~((mul_22_25_n_360 | mul_22_25_n_432) & (mul_22_25_n_615 | mul_22_25_n_433));
 assign mul_22_25_n_989 = ~((mul_22_25_n_354 | mul_22_25_n_279) & (mul_22_25_n_612 | mul_22_25_n_327));
 assign mul_22_25_n_988 = ~((mul_22_25_n_352 | mul_22_25_n_423) & (mul_22_25_n_604 | mul_22_25_n_237));
 assign mul_22_25_n_987 = ~((mul_22_25_n_355 | mul_22_25_n_99) & (mul_22_25_n_598 | mul_22_25_n_276));
 assign mul_22_25_n_986 = ~((mul_22_25_n_358 | mul_22_25_n_218) & (mul_22_25_n_613 | mul_22_25_n_210));
 assign mul_22_25_n_985 = ~((mul_22_25_n_358 | mul_22_25_n_509) & (mul_22_25_n_613 | mul_22_25_n_510));
 assign mul_22_25_n_984 = ~((mul_22_25_n_361 | mul_22_25_n_158) & (mul_22_25_n_616 | mul_22_25_n_142));
 assign mul_22_25_n_983 = ~((mul_22_25_n_350 | mul_22_25_n_467) & (mul_22_25_n_606 | mul_22_25_n_478));
 assign mul_22_25_n_982 = ~((mul_22_25_n_356 | mul_22_25_n_252) & (mul_22_25_n_600 | mul_22_25_n_416));
 assign mul_22_25_n_981 = ~((mul_22_25_n_352 | mul_22_25_n_247) & (mul_22_25_n_604 | mul_22_25_n_306));
 assign mul_22_25_n_980 = ~((mul_22_25_n_358 | mul_22_25_n_219) & (mul_22_25_n_613 | mul_22_25_n_213));
 assign mul_22_25_n_979 = ~((mul_22_25_n_363 | mul_22_25_n_120) & (mul_22_25_n_618 | mul_22_25_n_111));
 assign mul_22_25_n_978 = ~((mul_22_25_n_351 | mul_22_25_n_516) & (mul_22_25_n_596 | mul_22_25_n_528));
 assign mul_22_25_n_977 = ~((mul_22_25_n_361 | mul_22_25_n_429) & (mul_22_25_n_616 | mul_22_25_n_183));
 assign mul_22_25_n_976 = ~((mul_22_25_n_350 | mul_22_25_n_245) & (mul_22_25_n_606 | mul_22_25_n_308));
 assign mul_22_25_n_975 = ~((mul_22_25_n_362 | mul_22_25_n_161) & (mul_22_25_n_617 | mul_22_25_n_137));
 assign mul_22_25_n_974 = ~((mul_22_25_n_349 | mul_22_25_n_571) & (mul_22_25_n_602 | mul_22_25_n_415));
 assign mul_22_25_n_973 = ~((mul_22_25_n_357 | mul_22_25_n_505) & (mul_22_25_n_608 | mul_22_25_n_506));
 assign mul_22_25_n_972 = ~((mul_22_25_n_363 | mul_22_25_n_107) & (mul_22_25_n_618 | mul_22_25_n_121));
 assign mul_22_25_n_971 = ~((mul_22_25_n_353 | mul_22_25_n_464) & (mul_22_25_n_610 | mul_22_25_n_476));
 assign mul_22_25_n_970 = ~((mul_22_25_n_352 | mul_22_25_n_227) & (mul_22_25_n_604 | mul_22_25_n_228));
 assign mul_22_25_n_969 = ~((mul_22_25_n_352 | mul_22_25_n_369) & (mul_22_25_n_604 | mul_22_25_n_398));
 assign mul_22_25_n_968 = ~((mul_22_25_n_352 | mul_22_25_n_502) & (mul_22_25_n_604 | mul_22_25_n_488));
 assign mul_22_25_n_967 = ~((mul_22_25_n_357 | mul_22_25_n_280) & (mul_22_25_n_608 | mul_22_25_n_324));
 assign mul_22_25_n_966 = ~((mul_22_25_n_349 | mul_22_25_n_447) & (mul_22_25_n_602 | mul_22_25_n_445));
 assign mul_22_25_n_965 = ~((mul_22_25_n_350 | mul_22_25_n_308) & (mul_22_25_n_606 | mul_22_25_n_410));
 assign mul_22_25_n_964 = ~((mul_22_25_n_360 | mul_22_25_n_433) & (mul_22_25_n_615 | mul_22_25_n_222));
 assign mul_22_25_n_963 = ~((mul_22_25_n_360 | mul_22_25_n_174) & (mul_22_25_n_615 | mul_22_25_n_180));
 assign mul_22_25_n_962 = ~((mul_22_25_n_352 | mul_22_25_n_387) & (mul_22_25_n_604 | mul_22_25_n_423));
 assign mul_22_25_n_961 = ~((mul_22_25_n_356 | mul_22_25_n_438) & (mul_22_25_n_600 | mul_22_25_n_439));
 assign mul_22_25_n_960 = ~((mul_22_25_n_353 | mul_22_25_n_385) & (mul_22_25_n_610 | mul_22_25_n_579));
 assign mul_22_25_n_959 = ~((mul_22_25_n_358 | mul_22_25_n_211) & (mul_22_25_n_613 | mul_22_25_n_207));
 assign mul_22_25_n_958 = ~((mul_22_25_n_357 | mul_22_25_n_328) & (mul_22_25_n_608 | mul_22_25_n_315));
 assign mul_22_25_n_957 = ~((mul_22_25_n_363 | mul_22_25_n_113) & (mul_22_25_n_618 | mul_22_25_n_117));
 assign mul_22_25_n_956 = ~((mul_22_25_n_354 | mul_22_25_n_322) & (mul_22_25_n_612 | mul_22_25_n_233));
 assign mul_22_25_n_955 = ~((mul_22_25_n_363 | mul_22_25_n_103) & (mul_22_25_n_618 | mul_22_25_n_118));
 assign mul_22_25_n_954 = ~((mul_22_25_n_358 | mul_22_25_n_458) & (mul_22_25_n_613 | mul_22_25_n_430));
 assign mul_22_25_n_953 = ~((mul_22_25_n_355 | mul_22_25_n_323) & (mul_22_25_n_598 | mul_22_25_n_413));
 assign mul_22_25_n_952 = ~((mul_22_25_n_362 | mul_22_25_n_135) & (mul_22_25_n_617 | mul_22_25_n_139));
 assign mul_22_25_n_951 = ~((mul_22_25_n_362 | mul_22_25_n_137) & (mul_22_25_n_617 | mul_22_25_n_130));
 assign mul_22_25_n_950 = ~((mul_22_25_n_352 | mul_22_25_n_288) & (mul_22_25_n_604 | mul_22_25_n_247));
 assign mul_22_25_n_949 = ~((mul_22_25_n_358 | mul_22_25_n_486) & (mul_22_25_n_613 | mul_22_25_n_459));
 assign mul_22_25_n_948 = ~((mul_22_25_n_349 | mul_22_25_n_500) & (mul_22_25_n_602 | mul_22_25_n_473));
 assign mul_22_25_n_947 = ~((mul_22_25_n_351 | mul_22_25_n_542) & (mul_22_25_n_596 | mul_22_25_n_516));
 assign mul_22_25_n_946 = ~((mul_22_25_n_355 | mul_22_25_n_372) & (mul_22_25_n_598 | mul_22_25_n_99));
 assign mul_22_25_n_945 = ~((mul_22_25_n_350 | mul_22_25_n_370) & (mul_22_25_n_606 | mul_22_25_n_245));
 assign mul_22_25_n_944 = ~((mul_22_25_n_353 | mul_22_25_n_388) & (mul_22_25_n_610 | mul_22_25_n_265));
 assign mul_22_25_n_943 = ~((mul_22_25_n_356 | mul_22_25_n_466) & (mul_22_25_n_600 | mul_22_25_n_438));
 assign mul_22_25_n_942 = ~((mul_22_25_n_350 | mul_22_25_n_424) & (mul_22_25_n_606 | mul_22_25_n_297));
 assign mul_22_25_n_941 = ~((mul_22_25_n_358 | mul_22_25_n_216) & (mul_22_25_n_613 | mul_22_25_n_220));
 assign mul_22_25_n_940 = ~((mul_22_25_n_352 | mul_22_25_n_521) & (mul_22_25_n_604 | mul_22_25_n_502));
 assign mul_22_25_n_939 = ~((mul_22_25_n_351 | mul_22_25_n_368) & (mul_22_25_n_596 | mul_22_25_n_286));
 assign mul_22_25_n_938 = ~((mul_22_25_n_351 | mul_22_25_n_532) & (mul_22_25_n_596 | mul_22_25_n_96));
 assign mul_22_25_n_937 = ~((mul_22_25_n_357 | mul_22_25_n_443) & (mul_22_25_n_608 | mul_22_25_n_404));
 assign mul_22_25_n_936 = ~((mul_22_25_n_359 | mul_22_25_n_192) & (mul_22_25_n_614 | mul_22_25_n_195));
 assign mul_22_25_n_935 = ~((mul_22_25_n_354 | mul_22_25_n_474) & (mul_22_25_n_612 | mul_22_25_n_452));
 assign mul_22_25_n_934 = ~((mul_22_25_n_355 | mul_22_25_n_401) & (mul_22_25_n_598 | mul_22_25_n_323));
 assign mul_22_25_n_933 = ~((mul_22_25_n_357 | mul_22_25_n_511) & (mul_22_25_n_608 | mul_22_25_n_505));
 assign mul_22_25_n_932 = ~((mul_22_25_n_354 | mul_22_25_n_231) & (mul_22_25_n_612 | mul_22_25_n_290));
 assign mul_22_25_n_931 = ~((mul_22_25_n_361 | mul_22_25_n_155) & (mul_22_25_n_616 | mul_22_25_n_150));
 assign mul_22_25_n_930 = ~((mul_22_25_n_356 | mul_22_25_n_296) & (mul_22_25_n_600 | mul_22_25_n_409));
 assign mul_22_25_n_929 = ~((mul_22_25_n_362 | mul_22_25_n_124) & (mul_22_25_n_617 | mul_22_25_n_132));
 assign mul_22_25_n_928 = ~((mul_22_25_n_350 | mul_22_25_n_297) & (mul_22_25_n_606 | mul_22_25_n_389));
 assign mul_22_25_n_927 = ~((mul_22_25_n_349 | mul_22_25_n_556) & (mul_22_25_n_602 | mul_22_25_n_529));
 assign mul_22_25_n_926 = ~((mul_22_25_n_362 | mul_22_25_n_125) & (mul_22_25_n_617 | mul_22_25_n_127));
 assign mul_22_25_n_925 = ~((mul_22_25_n_358 | mul_22_25_n_212) & (mul_22_25_n_613 | mul_22_25_n_203));
 assign mul_22_25_n_924 = ~((mul_22_25_n_357 | mul_22_25_n_375) & (mul_22_25_n_608 | mul_22_25_n_280));
 assign mul_22_25_n_923 = ~((mul_22_25_n_356 | mul_22_25_n_311) & (mul_22_25_n_600 | mul_22_25_n_95));
 assign mul_22_25_n_922 = ~((mul_22_25_n_349 | mul_22_25_n_580) & (mul_22_25_n_602 | mul_22_25_n_364));
 assign mul_22_25_n_921 = ~((mul_22_25_n_361 | mul_22_25_n_183) & (mul_22_25_n_616 | mul_22_25_n_182));
 assign mul_22_25_n_920 = ~((mul_22_25_n_349 | mul_22_25_n_326) & (mul_22_25_n_602 | mul_22_25_n_580));
 assign mul_22_25_n_919 = ~((mul_22_25_n_353 | mul_22_25_n_497) & (mul_22_25_n_610 | mul_22_25_n_464));
 assign mul_22_25_n_918 = ~((mul_22_25_n_351 | mul_22_25_n_379) & (mul_22_25_n_596 | mul_22_25_n_100));
 assign mul_22_25_n_917 = ~((mul_22_25_n_357 | mul_22_25_n_325) & (mul_22_25_n_608 | mul_22_25_n_281));
 assign mul_22_25_n_1143 = ~(mul_22_25_n_664 & mul_22_25_n_637);
 assign mul_22_25_n_1142 = ~((mul_22_25_n_351 | mul_22_25_n_585) & (mul_22_25_n_596 | mul_22_25_n_72));
 assign mul_22_25_n_1139 = ~(mul_22_25_n_619 | (mul_22_25_n_595 & mul_22_25_n_576));
 assign mul_22_25_n_1137 = ~(mul_22_25_n_3 & (mul_22_25_n_606 | mul_22_25_n_562));
 assign mul_22_25_n_1134 = ~((mul_22_25_n_593 & mul_22_25_n_552) | (mul_22_25_n_601 & mul_22_25_n_557));
 assign mul_22_25_n_1133 = ~(mul_22_25_n_664 | mul_22_25_n_637);
 assign mul_22_25_n_1132 = ~((mul_22_25_n_594 & mul_22_25_n_472) | (mul_22_25_n_595 & mul_22_25_n_470));
 assign mul_22_25_n_1131 = ~((mul_22_25_n_351 | mul_22_25_n_286) & (mul_22_25_n_596 | mul_22_25_n_284));
 assign mul_22_25_n_1130 = ~(mul_22_25_n_679 & {in2[15]});
 assign mul_22_25_n_1129 = ~(mul_22_25_n_667 & {in2[17]});
 assign mul_22_25_n_1128 = ~(mul_22_25_n_680 & {in2[9]});
 assign mul_22_25_n_1127 = ~(mul_22_25_n_669 & {in2[5]});
 assign mul_22_25_n_1126 = ~(mul_22_25_n_671 & {in2[13]});
 assign mul_22_25_n_1125 = ~(mul_22_25_n_675 & {in2[7]});
 assign mul_22_25_n_1124 = ~(mul_22_25_n_676 & {in2[11]});
 assign mul_22_25_n_1123 = ~(mul_22_25_n_678 & {in2[19]});
 assign mul_22_25_n_1122 = ~(mul_22_25_n_681 & {in2[3]});
 assign mul_22_25_n_1121 = ~(mul_22_25_n_673 & {in2[21]});
 assign mul_22_25_n_1120 = ~(mul_22_25_n_672 & {in2[23]});
 assign mul_22_25_n_1119 = ~(mul_22_25_n_670 & {in2[25]});
 assign mul_22_25_n_1118 = ~(mul_22_25_n_668 & {in2[27]});
 assign mul_22_25_n_1117 = ~(mul_22_25_n_677 & {in2[29]});
 assign mul_22_25_n_1116 = ~(mul_22_25_n_674 & {in2[31]});
 assign mul_22_25_n_1115 = ~((mul_22_25_n_594 & mul_22_25_n_406) | (mul_22_25_n_595 & mul_22_25_n_428));
 assign mul_22_25_n_1114 = ~((mul_22_25_n_351 | mul_22_25_n_403) & (mul_22_25_n_596 | mul_22_25_n_532));
 assign mul_22_25_n_1113 = ~(mul_22_25_n_687 | mul_22_25_n_508);
 assign mul_22_25_n_916 = ~mul_22_25_n_915;
 assign mul_22_25_n_913 = ~mul_22_25_n_912;
 assign mul_22_25_n_911 = ~mul_22_25_n_910;
 assign mul_22_25_n_907 = ~((mul_22_25_n_356 | mul_22_25_n_160) & (mul_22_25_n_600 | mul_22_25_n_278));
 assign mul_22_25_n_906 = ~((mul_22_25_n_351 | mul_22_25_n_391) & (mul_22_25_n_596 | mul_22_25_n_282));
 assign mul_22_25_n_905 = ~((mul_22_25_n_349 | mul_22_25_n_364) & (mul_22_25_n_602 | mul_22_25_n_258));
 assign mul_22_25_n_904 = ~((mul_22_25_n_359 | mul_22_25_n_191) & (mul_22_25_n_614 | mul_22_25_n_189));
 assign mul_22_25_n_903 = ~((mul_22_25_n_352 | mul_22_25_n_312) & (mul_22_25_n_604 | mul_22_25_n_254));
 assign mul_22_25_n_902 = ~((mul_22_25_n_355 | mul_22_25_n_314) & (mul_22_25_n_598 | mul_22_25_n_401));
 assign mul_22_25_n_901 = ~((mul_22_25_n_360 | mul_22_25_n_169) & (mul_22_25_n_615 | mul_22_25_n_164));
 assign mul_22_25_n_900 = ~((mul_22_25_n_351 | mul_22_25_n_528) & (mul_22_25_n_596 | mul_22_25_n_490));
 assign mul_22_25_n_899 = ~((mul_22_25_n_357 | mul_22_25_n_94) & (mul_22_25_n_608 | mul_22_25_n_375));
 assign mul_22_25_n_898 = ~((mul_22_25_n_358 | mul_22_25_n_459) & (mul_22_25_n_613 | mul_22_25_n_458));
 assign mul_22_25_n_897 = ~((mul_22_25_n_356 | mul_22_25_n_287) & (mul_22_25_n_600 | mul_22_25_n_311));
 assign mul_22_25_n_896 = ~((mul_22_25_n_351 | mul_22_25_n_96) & (mul_22_25_n_596 | mul_22_25_n_181));
 assign mul_22_25_n_895 = ~((mul_22_25_n_355 | mul_22_25_n_525) & (mul_22_25_n_598 | mul_22_25_n_496));
 assign mul_22_25_n_894 = ~((mul_22_25_n_363 | mul_22_25_n_106) & (mul_22_25_n_618 | mul_22_25_n_108));
 assign mul_22_25_n_893 = ~((mul_22_25_n_350 | mul_22_25_n_587) & (mul_22_25_n_606 | mul_22_25_n_272));
 assign mul_22_25_n_892 = ~((mul_22_25_n_356 | mul_22_25_n_493) & (mul_22_25_n_600 | mul_22_25_n_477));
 assign mul_22_25_n_891 = ~((mul_22_25_n_354 | mul_22_25_n_588) & (mul_22_25_n_612 | mul_22_25_n_318));
 assign mul_22_25_n_890 = ~((mul_22_25_n_352 | mul_22_25_n_306) & (mul_22_25_n_604 | mul_22_25_n_384));
 assign mul_22_25_n_889 = ~((mul_22_25_n_358 | mul_22_25_n_217) & (mul_22_25_n_613 | mul_22_25_n_215));
 assign mul_22_25_n_888 = ~((mul_22_25_n_353 | mul_22_25_n_377) & (mul_22_25_n_610 | mul_22_25_n_321));
 assign mul_22_25_n_887 = ~((mul_22_25_n_352 | mul_22_25_n_543) & (mul_22_25_n_604 | mul_22_25_n_512));
 assign mul_22_25_n_886 = ~((mul_22_25_n_357 | mul_22_25_n_422) & (mul_22_25_n_608 | mul_22_25_n_325));
 assign mul_22_25_n_885 = ~((mul_22_25_n_357 | mul_22_25_n_482) & (mul_22_25_n_608 | mul_22_25_n_455));
 assign mul_22_25_n_884 = ~((mul_22_25_n_358 | mul_22_25_n_531) & (mul_22_25_n_613 | mul_22_25_n_509));
 assign mul_22_25_n_883 = ~((mul_22_25_n_352 | mul_22_25_n_555) & (mul_22_25_n_604 | mul_22_25_n_543));
 assign mul_22_25_n_882 = ~((mul_22_25_n_359 | mul_22_25_n_198) & (mul_22_25_n_614 | mul_22_25_n_202));
 assign mul_22_25_n_881 = ~((mul_22_25_n_360 | mul_22_25_n_172) & (mul_22_25_n_615 | mul_22_25_n_179));
 assign mul_22_25_n_880 = ~((mul_22_25_n_349 | mul_22_25_n_445) & (mul_22_25_n_602 | mul_22_25_n_263));
 assign mul_22_25_n_879 = ~((mul_22_25_n_351 | mul_22_25_n_282) & (mul_22_25_n_596 | mul_22_25_n_585));
 assign mul_22_25_n_878 = ~((mul_22_25_n_361 | mul_22_25_n_144) & (mul_22_25_n_616 | mul_22_25_n_143));
 assign mul_22_25_n_877 = ~((mul_22_25_n_362 | mul_22_25_n_131) & (mul_22_25_n_617 | mul_22_25_n_134));
 assign mul_22_25_n_876 = ~((mul_22_25_n_352 | mul_22_25_n_488) & (mul_22_25_n_604 | mul_22_25_n_462));
 assign mul_22_25_n_875 = ~((mul_22_25_n_353 | mul_22_25_n_394) & (mul_22_25_n_610 | mul_22_25_n_383));
 assign mul_22_25_n_874 = ~((mul_22_25_n_355 | mul_22_25_n_503) & (mul_22_25_n_598 | mul_22_25_n_481));
 assign mul_22_25_n_873 = ~((mul_22_25_n_353 | mul_22_25_n_553) & (mul_22_25_n_610 | mul_22_25_n_534));
 assign mul_22_25_n_872 = ~((mul_22_25_n_354 | mul_22_25_n_452) & (mul_22_25_n_612 | mul_22_25_n_451));
 assign mul_22_25_n_871 = ~((mul_22_25_n_353 | mul_22_25_n_91) & (mul_22_25_n_610 | mul_22_25_n_395));
 assign mul_22_25_n_870 = ~((mul_22_25_n_357 | mul_22_25_n_378) & (mul_22_25_n_608 | mul_22_25_n_238));
 assign mul_22_25_n_869 = ~((mul_22_25_n_356 | mul_22_25_n_581) & (mul_22_25_n_600 | mul_22_25_n_371));
 assign mul_22_25_n_868 = ~((mul_22_25_n_350 | mul_22_25_n_487) & (mul_22_25_n_606 | mul_22_25_n_492));
 assign mul_22_25_n_867 = ~((mul_22_25_n_351 | mul_22_25_n_444) & (mul_22_25_n_596 | mul_22_25_n_403));
 assign mul_22_25_n_866 = ~((mul_22_25_n_357 | mul_22_25_n_295) & (mul_22_25_n_608 | mul_22_25_n_98));
 assign mul_22_25_n_865 = ~((mul_22_25_n_350 | mul_22_25_n_101) & (mul_22_25_n_606 | mul_22_25_n_367));
 assign mul_22_25_n_864 = ~((mul_22_25_n_355 | mul_22_25_n_300) & (mul_22_25_n_598 | mul_22_25_n_460));
 assign mul_22_25_n_863 = ~((mul_22_25_n_355 | mul_22_25_n_481) & (mul_22_25_n_598 | mul_22_25_n_480));
 assign mul_22_25_n_862 = ~((mul_22_25_n_358 | mul_22_25_n_430) & (mul_22_25_n_613 | mul_22_25_n_431));
 assign mul_22_25_n_861 = ~((mul_22_25_n_349 | mul_22_25_n_258) & (mul_22_25_n_602 | mul_22_25_n_400));
 assign mul_22_25_n_860 = ~((mul_22_25_n_354 | mul_22_25_n_537) & (mul_22_25_n_612 | mul_22_25_n_548));
 assign mul_22_25_n_859 = ~((mul_22_25_n_350 | mul_22_25_n_88) & (mul_22_25_n_606 | mul_22_25_n_285));
 assign mul_22_25_n_858 = ~((mul_22_25_n_356 | mul_22_25_n_402) & (mul_22_25_n_600 | mul_22_25_n_242));
 assign mul_22_25_n_857 = ~((mul_22_25_n_356 | mul_22_25_n_495) & (mul_22_25_n_600 | mul_22_25_n_493));
 assign mul_22_25_n_856 = ~((mul_22_25_n_353 | mul_22_25_n_86) & (mul_22_25_n_610 | mul_22_25_n_385));
 assign mul_22_25_n_855 = ~((mul_22_25_n_360 | mul_22_25_n_170) & (mul_22_25_n_615 | mul_22_25_n_166));
 assign mul_22_25_n_854 = ~((mul_22_25_n_354 | mul_22_25_n_421) & (mul_22_25_n_612 | mul_22_25_n_366));
 assign mul_22_25_n_853 = ~((mul_22_25_n_357 | mul_22_25_n_475) & (mul_22_25_n_608 | mul_22_25_n_482));
 assign mul_22_25_n_852 = ~((mul_22_25_n_358 | mul_22_25_n_214) & (mul_22_25_n_613 | mul_22_25_n_217));
 assign mul_22_25_n_851 = ~((mul_22_25_n_359 | mul_22_25_n_193) & (mul_22_25_n_614 | mul_22_25_n_198));
 assign mul_22_25_n_850 = ~((mul_22_25_n_355 | mul_22_25_n_524) & (mul_22_25_n_598 | mul_22_25_n_525));
 assign mul_22_25_n_849 = ~((mul_22_25_n_352 | mul_22_25_n_97) & (mul_22_25_n_604 | mul_22_25_n_312));
 assign mul_22_25_n_848 = ~((mul_22_25_n_361 | mul_22_25_n_147) & (mul_22_25_n_616 | mul_22_25_n_144));
 assign mul_22_25_n_847 = ~((mul_22_25_n_350 | mul_22_25_n_273) & (mul_22_25_n_606 | mul_22_25_n_587));
 assign mul_22_25_n_846 = ~((mul_22_25_n_356 | mul_22_25_n_95) & (mul_22_25_n_600 | mul_22_25_n_581));
 assign mul_22_25_n_845 = ~((mul_22_25_n_351 | mul_22_25_n_365) & (mul_22_25_n_596 | mul_22_25_n_275));
 assign mul_22_25_n_844 = ~((mul_22_25_n_357 | mul_22_25_n_405) & (mul_22_25_n_608 | mul_22_25_n_94));
 assign mul_22_25_n_843 = ~((mul_22_25_n_349 | mul_22_25_n_102) & (mul_22_25_n_602 | mul_22_25_n_326));
 assign mul_22_25_n_842 = ~((mul_22_25_n_363 | mul_22_25_n_105) & (mul_22_25_n_618 | mul_22_25_n_106));
 assign mul_22_25_n_841 = ~((mul_22_25_n_351 | mul_22_25_n_275) & (mul_22_25_n_596 | mul_22_25_n_303));
 assign mul_22_25_n_840 = ~((mul_22_25_n_354 | mul_22_25_n_327) & (mul_22_25_n_612 | mul_22_25_n_322));
 assign mul_22_25_n_839 = ~((mul_22_25_n_359 | mul_22_25_n_190) & (mul_22_25_n_614 | mul_22_25_n_199));
 assign mul_22_25_n_838 = ~(mul_22_25_n_684 & (mul_22_25_n_351 | mul_22_25_n_284));
 assign mul_22_25_n_837 = ~((mul_22_25_n_352 | mul_22_25_n_268) & (mul_22_25_n_604 | mul_22_25_n_97));
 assign mul_22_25_n_836 = ~((mul_22_25_n_363 | mul_22_25_n_104) & (mul_22_25_n_618 | mul_22_25_n_112));
 assign mul_22_25_n_835 = ~((mul_22_25_n_353 | mul_22_25_n_321) & (mul_22_25_n_610 | mul_22_25_n_411));
 assign mul_22_25_n_834 = ~((mul_22_25_n_353 | mul_22_25_n_453) & (mul_22_25_n_610 | mul_22_25_n_390));
 assign mul_22_25_n_833 = ~((mul_22_25_n_355 | mul_22_25_n_276) & (mul_22_25_n_598 | mul_22_25_n_381));
 assign mul_22_25_n_832 = ~((mul_22_25_n_355 | mul_22_25_n_584) & (mul_22_25_n_598 | mul_22_25_n_314));
 assign mul_22_25_n_831 = ~((mul_22_25_n_359 | mul_22_25_n_457) & (mul_22_25_n_614 | mul_22_25_n_426));
 assign mul_22_25_n_830 = ~((mul_22_25_n_361 | mul_22_25_n_159) & (mul_22_25_n_616 | mul_22_25_n_145));
 assign mul_22_25_n_829 = ~((mul_22_25_n_355 | mul_22_25_n_89) & (mul_22_25_n_598 | mul_22_25_n_225));
 assign mul_22_25_n_828 = ~((mul_22_25_n_350 | mul_22_25_n_523) & (mul_22_25_n_606 | mul_22_25_n_518));
 assign mul_22_25_n_827 = ~((mul_22_25_n_356 | mul_22_25_n_313) & (mul_22_25_n_600 | mul_22_25_n_287));
 assign mul_22_25_n_826 = ((mul_22_25_n_592 & mul_22_25_n_577) | (mul_22_25_n_611 & mul_22_25_n_538));
 assign mul_22_25_n_825 = ~((mul_22_25_n_356 | mul_22_25_n_302) & (mul_22_25_n_600 | mul_22_25_n_252));
 assign mul_22_25_n_824 = ~((mul_22_25_n_352 | mul_22_25_n_558) & (mul_22_25_n_604 | mul_22_25_n_555));
 assign mul_22_25_n_823 = ~((mul_22_25_n_350 | mul_22_25_n_540) & (mul_22_25_n_606 | mul_22_25_n_541));
 assign mul_22_25_n_822 = ~((mul_22_25_n_356 | mul_22_25_n_519) & (mul_22_25_n_600 | mul_22_25_n_495));
 assign mul_22_25_n_821 = ~((mul_22_25_n_353 | mul_22_25_n_248) & (mul_22_25_n_610 | mul_22_25_n_86));
 assign mul_22_25_n_820 = ~((mul_22_25_n_356 | mul_22_25_n_439) & (mul_22_25_n_600 | mul_22_25_n_386));
 assign mul_22_25_n_819 = ~((mul_22_25_n_354 | mul_22_25_n_309) & (mul_22_25_n_612 | mul_22_25_n_115));
 assign mul_22_25_n_818 = ~((mul_22_25_n_350 | mul_22_25_n_224) & (mul_22_25_n_606 | mul_22_25_n_88));
 assign mul_22_25_n_817 = ~((mul_22_25_n_355 | mul_22_25_n_533) & (mul_22_25_n_598 | mul_22_25_n_524));
 assign mul_22_25_n_816 = ~((mul_22_25_n_353 | mul_22_25_n_383) & (mul_22_25_n_610 | mul_22_25_n_91));
 assign mul_22_25_n_815 = ~((mul_22_25_n_355 | mul_22_25_n_436) & (mul_22_25_n_598 | mul_22_25_n_259));
 assign mul_22_25_n_814 = ~((mul_22_25_n_362 | mul_22_25_n_130) & (mul_22_25_n_617 | mul_22_25_n_133));
 assign mul_22_25_n_813 = ~((mul_22_25_n_357 | mul_22_25_n_238) & (mul_22_25_n_608 | mul_22_25_n_422));
 assign mul_22_25_n_812 = ~((mul_22_25_n_351 | mul_22_25_n_303) & (mul_22_25_n_596 | mul_22_25_n_368));
 assign mul_22_25_n_811 = ~((mul_22_25_n_360 | mul_22_25_n_167) & (mul_22_25_n_615 | mul_22_25_n_176));
 assign mul_22_25_n_810 = ~((mul_22_25_n_354 | mul_22_25_n_419) & (mul_22_25_n_612 | mul_22_25_n_421));
 assign mul_22_25_n_809 = ~((mul_22_25_n_350 | mul_22_25_n_440) & (mul_22_25_n_606 | mul_22_25_n_273));
 assign mul_22_25_n_808 = ~((mul_22_25_n_362 | mul_22_25_n_123) & (mul_22_25_n_617 | mul_22_25_n_138));
 assign mul_22_25_n_807 = ~((mul_22_25_n_363 | mul_22_25_n_112) & (mul_22_25_n_618 | mul_22_25_n_105));
 assign mul_22_25_n_806 = ~((mul_22_25_n_358 | mul_22_25_n_206) & (mul_22_25_n_613 | mul_22_25_n_211));
 assign mul_22_25_n_805 = ~((mul_22_25_n_362 | mul_22_25_n_127) & (mul_22_25_n_617 | mul_22_25_n_126));
 assign mul_22_25_n_804 = ~((mul_22_25_n_359 | mul_22_25_n_484) & (mul_22_25_n_614 | mul_22_25_n_456));
 assign mul_22_25_n_803 = ~((mul_22_25_n_349 | mul_22_25_n_396) & (mul_22_25_n_602 | mul_22_25_n_102));
 assign mul_22_25_n_802 = ~((mul_22_25_n_354 | mul_22_25_n_289) & (mul_22_25_n_612 | mul_22_25_n_309));
 assign mul_22_25_n_801 = ~((mul_22_25_n_350 | mul_22_25_n_389) & (mul_22_25_n_606 | mul_22_25_n_380));
 assign mul_22_25_n_800 = ~((mul_22_25_n_358 | mul_22_25_n_205) & (mul_22_25_n_613 | mul_22_25_n_204));
 assign mul_22_25_n_799 = ~((mul_22_25_n_355 | mul_22_25_n_259) & (mul_22_25_n_598 | mul_22_25_n_420));
 assign mul_22_25_n_798 = ~((mul_22_25_n_363 | mul_22_25_n_121) & (mul_22_25_n_618 | mul_22_25_n_119));
 assign mul_22_25_n_797 = ~((mul_22_25_n_350 | mul_22_25_n_446) & (mul_22_25_n_606 | mul_22_25_n_440));
 assign mul_22_25_n_796 = ~((mul_22_25_n_361 | mul_22_25_n_153) & (mul_22_25_n_616 | mul_22_25_n_148));
 assign mul_22_25_n_795 = ~((mul_22_25_n_357 | mul_22_25_n_569) & (mul_22_25_n_608 | mul_22_25_n_535));
 assign mul_22_25_n_794 = ~((mul_22_25_n_353 | mul_22_25_n_390) & (mul_22_25_n_610 | mul_22_25_n_248));
 assign mul_22_25_n_793 = ~((mul_22_25_n_363 | mul_22_25_n_119) & (mul_22_25_n_618 | mul_22_25_n_110));
 assign mul_22_25_n_792 = ~((mul_22_25_n_351 | mul_22_25_n_274) & (mul_22_25_n_596 | mul_22_25_n_391));
 assign mul_22_25_n_791 = ~((mul_22_25_n_355 | mul_22_25_n_226) & (mul_22_25_n_598 | mul_22_25_n_584));
 assign mul_22_25_n_790 = ~((mul_22_25_n_354 | mul_22_25_n_465) & (mul_22_25_n_612 | mul_22_25_n_474));
 assign mul_22_25_n_789 = ~((mul_22_25_n_354 | mul_22_25_n_283) & (mul_22_25_n_612 | mul_22_25_n_373));
 assign mul_22_25_n_788 = ~((mul_22_25_n_353 | mul_22_25_n_319) & (mul_22_25_n_610 | mul_22_25_n_307));
 assign mul_22_25_n_787 = ((mul_22_25_n_594 & mul_22_25_n_470) | (mul_22_25_n_595 & mul_22_25_n_449));
 assign mul_22_25_n_786 = ~((mul_22_25_n_356 | mul_22_25_n_264) & (mul_22_25_n_600 | mul_22_25_n_313));
 assign mul_22_25_n_785 = ~((mul_22_25_n_355 | mul_22_25_n_420) & (mul_22_25_n_598 | mul_22_25_n_87));
 assign mul_22_25_n_784 = ~((mul_22_25_n_357 | mul_22_25_n_324) & (mul_22_25_n_608 | mul_22_25_n_295));
 assign mul_22_25_n_783 = ~((mul_22_25_n_357 | mul_22_25_n_315) & (mul_22_25_n_608 | mul_22_25_n_262));
 assign mul_22_25_n_782 = ~((mul_22_25_n_358 | mul_22_25_n_208) & (mul_22_25_n_613 | mul_22_25_n_209));
 assign mul_22_25_n_781 = ~((mul_22_25_n_355 | mul_22_25_n_564) & (mul_22_25_n_598 | mul_22_25_n_539));
 assign mul_22_25_n_780 = ~((mul_22_25_n_350 | mul_22_25_n_367) & (mul_22_25_n_606 | mul_22_25_n_224));
 assign mul_22_25_n_779 = ~((mul_22_25_n_351 | mul_22_25_n_239) & (mul_22_25_n_596 | mul_22_25_n_274));
 assign mul_22_25_n_778 = ~((mul_22_25_n_354 | mul_22_25_n_373) & (mul_22_25_n_612 | mul_22_25_n_289));
 assign mul_22_25_n_777 = ~((mul_22_25_n_358 | mul_22_25_n_210) & (mul_22_25_n_613 | mul_22_25_n_205));
 assign mul_22_25_n_776 = ~((mul_22_25_n_356 | mul_22_25_n_416) & (mul_22_25_n_600 | mul_22_25_n_257));
 assign mul_22_25_n_775 = ~((mul_22_25_n_360 | mul_22_25_n_163) & (mul_22_25_n_615 | mul_22_25_n_178));
 assign mul_22_25_n_774 = ~((mul_22_25_n_354 | mul_22_25_n_253) & (mul_22_25_n_612 | mul_22_25_n_419));
 assign mul_22_25_n_773 = ~((mul_22_25_n_352 | mul_22_25_n_392) & (mul_22_25_n_604 | mul_22_25_n_414));
 assign mul_22_25_n_772 = ~((mul_22_25_n_350 | mul_22_25_n_478) & (mul_22_25_n_606 | mul_22_25_n_446));
 assign mul_22_25_n_771 = ~((mul_22_25_n_349 | mul_22_25_n_269) & (mul_22_25_n_602 | mul_22_25_n_271));
 assign mul_22_25_n_770 = ~((mul_22_25_n_361 | mul_22_25_n_152) & (mul_22_25_n_616 | mul_22_25_n_153));
 assign mul_22_25_n_769 = ~((mul_22_25_n_362 | mul_22_25_n_136) & (mul_22_25_n_617 | mul_22_25_n_128));
 assign mul_22_25_n_768 = ~((mul_22_25_n_354 | mul_22_25_n_366) & (mul_22_25_n_612 | mul_22_25_n_231));
 assign mul_22_25_n_767 = ~((mul_22_25_n_362 | mul_22_25_n_128) & (mul_22_25_n_617 | mul_22_25_n_123));
 assign mul_22_25_n_766 = ~((mul_22_25_n_349 | mul_22_25_n_301) & (mul_22_25_n_602 | mul_22_25_n_396));
 assign mul_22_25_n_765 = ~((mul_22_25_n_357 | mul_22_25_n_404) & (mul_22_25_n_608 | mul_22_25_n_328));
 assign mul_22_25_n_764 = ~((mul_22_25_n_354 | mul_22_25_n_310) & (mul_22_25_n_612 | mul_22_25_n_279));
 assign mul_22_25_n_763 = ~((mul_22_25_n_350 | mul_22_25_n_562) & (mul_22_25_n_606 | mul_22_25_n_540));
 assign mul_22_25_n_762 = ~((mul_22_25_n_349 | mul_22_25_n_501) & (mul_22_25_n_602 | mul_22_25_n_500));
 assign mul_22_25_n_761 = ~((mul_22_25_n_360 | mul_22_25_n_177) & (mul_22_25_n_615 | mul_22_25_n_163));
 assign mul_22_25_n_760 = ~((mul_22_25_n_359 | mul_22_25_n_199) & (mul_22_25_n_614 | mul_22_25_n_186));
 assign mul_22_25_n_759 = ~((mul_22_25_n_363 | mul_22_25_n_118) & (mul_22_25_n_618 | mul_22_25_n_116));
 assign mul_22_25_n_758 = ~((mul_22_25_n_357 | mul_22_25_n_583) & (mul_22_25_n_608 | mul_22_25_n_578));
 assign mul_22_25_n_757 = ~((mul_22_25_n_362 | mul_22_25_n_140) & (mul_22_25_n_617 | mul_22_25_n_136));
 assign mul_22_25_n_756 = ~((mul_22_25_n_357 | mul_22_25_n_514) & (mul_22_25_n_608 | mul_22_25_n_511));
 assign mul_22_25_n_755 = ~((mul_22_25_n_358 | mul_22_25_n_203) & (mul_22_25_n_613 | mul_22_25_n_206));
 assign mul_22_25_n_754 = ~((mul_22_25_n_361 | mul_22_25_n_182) & (mul_22_25_n_616 | mul_22_25_n_159));
 assign mul_22_25_n_753 = ~((mul_22_25_n_352 | mul_22_25_n_237) & (mul_22_25_n_604 | mul_22_25_n_241));
 assign mul_22_25_n_752 = ~((mul_22_25_n_356 | mul_22_25_n_257) & (mul_22_25_n_600 | mul_22_25_n_402));
 assign mul_22_25_n_751 = ~((mul_22_25_n_354 | mul_22_25_n_499) & (mul_22_25_n_612 | mul_22_25_n_465));
 assign mul_22_25_n_750 = ~((mul_22_25_n_349 | mul_22_25_n_271) & (mul_22_25_n_602 | mul_22_25_n_230));
 assign mul_22_25_n_749 = ~((mul_22_25_n_351 | mul_22_25_n_100) & (mul_22_25_n_596 | mul_22_25_n_365));
 assign mul_22_25_n_748 = ~((mul_22_25_n_353 | mul_22_25_n_307) & (mul_22_25_n_610 | mul_22_25_n_394));
 assign mul_22_25_n_747 = ~((mul_22_25_n_355 | mul_22_25_n_413) & (mul_22_25_n_598 | mul_22_25_n_291));
 assign mul_22_25_n_746 = ~((mul_22_25_n_350 | mul_22_25_n_320) & (mul_22_25_n_606 | mul_22_25_n_101));
 assign mul_22_25_n_745 = ~((mul_22_25_n_360 | mul_22_25_n_162) & (mul_22_25_n_615 | mul_22_25_n_169));
 assign mul_22_25_n_744 = ~((mul_22_25_n_363 | mul_22_25_n_109) & (mul_22_25_n_618 | mul_22_25_n_113));
 assign mul_22_25_n_743 = ~((mul_22_25_n_360 | mul_22_25_n_180) & (mul_22_25_n_615 | mul_22_25_n_170));
 assign mul_22_25_n_742 = ~((mul_22_25_n_353 | mul_22_25_n_586) & (mul_22_25_n_610 | mul_22_25_n_412));
 assign mul_22_25_n_741 = ~((mul_22_25_n_356 | mul_22_25_n_574) & (mul_22_25_n_600 | mul_22_25_n_536));
 assign mul_22_25_n_740 = ~((mul_22_25_n_350 | mul_22_25_n_90) & (mul_22_25_n_606 | mul_22_25_n_266));
 assign mul_22_25_n_739 = ~((mul_22_25_n_358 | mul_22_25_n_209) & (mul_22_25_n_613 | mul_22_25_n_218));
 assign mul_22_25_n_738 = ~((mul_22_25_n_355 | mul_22_25_n_246) & (mul_22_25_n_598 | mul_22_25_n_226));
 assign mul_22_25_n_737 = ~((mul_22_25_n_359 | mul_22_25_n_189) & (mul_22_25_n_614 | mul_22_25_n_194));
 assign mul_22_25_n_736 = ~((mul_22_25_n_350 | mul_22_25_n_492) & (mul_22_25_n_606 | mul_22_25_n_467));
 assign mul_22_25_n_735 = ~((mul_22_25_n_357 | mul_22_25_n_229) & (mul_22_25_n_608 | mul_22_25_n_583));
 assign mul_22_25_n_734 = ~((mul_22_25_n_360 | mul_22_25_n_171) & (mul_22_25_n_615 | mul_22_25_n_177));
 assign mul_22_25_n_733 = ~((mul_22_25_n_359 | mul_22_25_n_186) & (mul_22_25_n_614 | mul_22_25_n_185));
 assign mul_22_25_n_732 = ~((mul_22_25_n_361 | mul_22_25_n_142) & (mul_22_25_n_616 | mul_22_25_n_154));
 assign mul_22_25_n_731 = ~((mul_22_25_n_357 | mul_22_25_n_544) & (mul_22_25_n_608 | mul_22_25_n_514));
 assign mul_22_25_n_730 = ~((mul_22_25_n_362 | mul_22_25_n_126) & (mul_22_25_n_617 | mul_22_25_n_140));
 assign mul_22_25_n_729 = ~((mul_22_25_n_352 | mul_22_25_n_254) & (mul_22_25_n_604 | mul_22_25_n_369));
 assign mul_22_25_n_728 = ~((mul_22_25_n_354 | mul_22_25_n_451) & (mul_22_25_n_612 | mul_22_25_n_283));
 assign mul_22_25_n_727 = ~((mul_22_25_n_353 | mul_22_25_n_448) & (mul_22_25_n_610 | mul_22_25_n_453));
 assign mul_22_25_n_726 = ~((mul_22_25_n_349 | mul_22_25_n_267) & (mul_22_25_n_602 | mul_22_25_n_269));
 assign mul_22_25_n_725 = ~((mul_22_25_n_359 | mul_22_25_n_185) & (mul_22_25_n_614 | mul_22_25_n_200));
 assign mul_22_25_n_724 = ~((mul_22_25_n_361 | mul_22_25_n_148) & (mul_22_25_n_616 | mul_22_25_n_147));
 assign mul_22_25_n_723 = ~((mul_22_25_n_352 | mul_22_25_n_241) & (mul_22_25_n_604 | mul_22_25_n_392));
 assign mul_22_25_n_722 = ~((mul_22_25_n_356 | mul_22_25_n_397) & (mul_22_25_n_600 | mul_22_25_n_264));
 assign mul_22_25_n_721 = ~((mul_22_25_n_356 | mul_22_25_n_242) & (mul_22_25_n_600 | mul_22_25_n_296));
 assign mul_22_25_n_720 = ~((mul_22_25_n_360 | mul_22_25_n_164) & (mul_22_25_n_615 | mul_22_25_n_171));
 assign mul_22_25_n_719 = ~((mul_22_25_n_349 | mul_22_25_n_463) & (mul_22_25_n_602 | mul_22_25_n_447));
 assign mul_22_25_n_718 = ~((mul_22_25_n_357 | mul_22_25_n_262) & (mul_22_25_n_608 | mul_22_25_n_229));
 assign mul_22_25_n_717 = ~((mul_22_25_n_360 | mul_22_25_n_165) & (mul_22_25_n_615 | mul_22_25_n_162));
 assign mul_22_25_n_716 = ~((mul_22_25_n_361 | mul_22_25_n_154) & (mul_22_25_n_616 | mul_22_25_n_152));
 assign mul_22_25_n_715 = ~((mul_22_25_n_358 | mul_22_25_n_204) & (mul_22_25_n_613 | mul_22_25_n_214));
 assign mul_22_25_n_714 = ((mul_22_25_n_594 & mul_22_25_n_428) | (mul_22_25_n_595 & mul_22_25_n_240));
 assign mul_22_25_n_713 = ~((mul_22_25_n_352 | mul_22_25_n_435) & (mul_22_25_n_604 | mul_22_25_n_268));
 assign mul_22_25_n_712 = ~((mul_22_25_n_359 | mul_22_25_n_195) & (mul_22_25_n_614 | mul_22_25_n_187));
 assign mul_22_25_n_711 = ~((mul_22_25_n_361 | mul_22_25_n_141) & (mul_22_25_n_616 | mul_22_25_n_149));
 assign mul_22_25_n_710 = ~((mul_22_25_n_361 | mul_22_25_n_143) & (mul_22_25_n_616 | mul_22_25_n_155));
 assign mul_22_25_n_709 = ~((mul_22_25_n_353 | mul_22_25_n_265) & (mul_22_25_n_610 | mul_22_25_n_586));
 assign mul_22_25_n_708 = ~((mul_22_25_n_359 | mul_22_25_n_507) & (mul_22_25_n_614 | mul_22_25_n_483));
 assign mul_22_25_n_707 = ~((mul_22_25_n_353 | mul_22_25_n_491) & (mul_22_25_n_610 | mul_22_25_n_497));
 assign mul_22_25_n_706 = ~((mul_22_25_n_350 | mul_22_25_n_410) & (mul_22_25_n_606 | mul_22_25_n_320));
 assign mul_22_25_n_705 = ~((mul_22_25_n_355 | mul_22_25_n_291) & (mul_22_25_n_598 | mul_22_25_n_89));
 assign mul_22_25_n_704 = ~((mul_22_25_n_355 | mul_22_25_n_381) & (mul_22_25_n_598 | mul_22_25_n_246));
 assign mul_22_25_n_703 = ~((mul_22_25_n_359 | mul_22_25_n_188) & (mul_22_25_n_614 | mul_22_25_n_191));
 assign mul_22_25_n_702 = ~((mul_22_25_n_350 | mul_22_25_n_380) & (mul_22_25_n_606 | mul_22_25_n_90));
 assign mul_22_25_n_701 = ~((mul_22_25_n_361 | mul_22_25_n_157) & (mul_22_25_n_616 | mul_22_25_n_158));
 assign mul_22_25_n_700 = ~((mul_22_25_n_349 | mul_22_25_n_374) & (mul_22_25_n_602 | mul_22_25_n_571));
 assign mul_22_25_n_699 = ~((mul_22_25_n_358 | mul_22_25_n_431) & (mul_22_25_n_613 | mul_22_25_n_208));
 assign mul_22_25_n_698 = ~((mul_22_25_n_363 | mul_22_25_n_116) & (mul_22_25_n_618 | mul_22_25_n_104));
 assign mul_22_25_n_697 = ~((mul_22_25_n_357 | mul_22_25_n_98) & (mul_22_25_n_608 | mul_22_25_n_378));
 assign mul_22_25_n_696 = ~((mul_22_25_n_352 | mul_22_25_n_469) & (mul_22_25_n_604 | mul_22_25_n_434));
 assign mul_22_25_n_695 = ~((mul_22_25_n_356 | mul_22_25_n_278) & (mul_22_25_n_600 | mul_22_25_n_397));
 assign mul_22_25_n_694 = ~((mul_22_25_n_357 | mul_22_25_n_578) & (mul_22_25_n_608 | mul_22_25_n_405));
 assign mul_22_25_n_693 = ~((mul_22_25_n_361 | mul_22_25_n_146) & (mul_22_25_n_616 | mul_22_25_n_157));
 assign mul_22_25_n_692 = ~((mul_22_25_n_360 | mul_22_25_n_175) & (mul_22_25_n_615 | mul_22_25_n_174));
 assign mul_22_25_n_691 = ~((mul_22_25_n_362 | mul_22_25_n_129) & (mul_22_25_n_617 | mul_22_25_n_125));
 assign mul_22_25_n_690 = ~((mul_22_25_n_359 | mul_22_25_n_196) & (mul_22_25_n_614 | mul_22_25_n_193));
 assign mul_22_25_n_689 = ~((mul_22_25_n_359 | mul_22_25_n_184) & (mul_22_25_n_614 | mul_22_25_n_188));
 assign mul_22_25_n_915 = ~((mul_22_25_n_356 | mul_22_25_n_536) & (mul_22_25_n_600 | mul_22_25_n_554));
 assign mul_22_25_n_914 = ~((~mul_22_25_n_596 & ~mul_22_25_n_545) | (mul_22_25_n_594 & mul_22_25_n_576));
 assign mul_22_25_n_912 = ~((mul_22_25_n_355 | mul_22_25_n_539) & (mul_22_25_n_598 | mul_22_25_n_533));
 assign mul_22_25_n_910 = ~((mul_22_25_n_357 | mul_22_25_n_535) & (mul_22_25_n_608 | mul_22_25_n_544));
 assign mul_22_25_n_909 = ((mul_22_25_n_351 | mul_22_25_n_490) & (mul_22_25_n_596 | mul_22_25_n_498));
 assign mul_22_25_n_908 = ~((mul_22_25_n_351 | mul_22_25_n_450) & (mul_22_25_n_596 | mul_22_25_n_444));
 assign mul_22_25_n_684 = ~(mul_22_25_n_595 & mul_22_25_n_406);
 assign mul_22_25_n_683 = ~((mul_22_25_n_504 | mul_22_25_n_26) & (mul_22_25_n_590 | mul_22_25_n_468));
 assign mul_22_25_n_682 = ~((mul_22_25_n_526 | mul_22_25_n_26) & (mul_22_25_n_590 | mul_22_25_n_527));
 assign mul_22_25_n_681 = ~(({in2[2]} & {in1[0]}) | ({in2[1]} & ({in2[2]} ^ {in1[0]})));
 assign mul_22_25_n_680 = ~(({in2[8]} & {in1[0]}) | ({in2[7]} & ({in2[8]} ^ {in1[0]})));
 assign mul_22_25_n_679 = ~(({in2[14]} & {in1[0]}) | ({in2[13]} & ({in2[14]} ^ {in1[0]})));
 assign mul_22_25_n_678 = ~(({in2[18]} & {in1[0]}) | ({in2[17]} & ({in2[18]} ^ {in1[0]})));
 assign mul_22_25_n_677 = ~(({in2[28]} & {in1[0]}) | ({in2[27]} & ({in2[28]} ^ {in1[0]})));
 assign mul_22_25_n_676 = ~(({in2[10]} & {in1[0]}) | ({in2[9]} & ({in2[10]} ^ {in1[0]})));
 assign mul_22_25_n_675 = ~(({in2[6]} & {in1[0]}) | ({in2[5]} & ({in2[6]} ^ {in1[0]})));
 assign mul_22_25_n_674 = ~(({in2[30]} & {in1[0]}) | ({in2[29]} & ({in2[30]} ^ {in1[0]})));
 assign mul_22_25_n_673 = ~(({in2[20]} & {in1[0]}) | ({in2[19]} & ({in2[20]} ^ {in1[0]})));
 assign mul_22_25_n_672 = ~(({in2[22]} & {in1[0]}) | ({in2[21]} & ({in2[22]} ^ {in1[0]})));
 assign mul_22_25_n_671 = ~(({in2[12]} & {in1[0]}) | ({in2[11]} & ({in2[12]} ^ {in1[0]})));
 assign mul_22_25_n_670 = ~(({in2[24]} & {in1[0]}) | ({in2[23]} & ({in2[24]} ^ {in1[0]})));
 assign mul_22_25_n_669 = ~(({in2[4]} & {in1[0]}) | ({in2[3]} & ({in2[4]} ^ {in1[0]})));
 assign mul_22_25_n_668 = ~(({in2[26]} & {in1[0]}) | ({in2[25]} & ({in2[26]} ^ {in1[0]})));
 assign mul_22_25_n_667 = ~(({in2[16]} & {in1[0]}) | ({in2[15]} & ({in2[16]} ^ {in1[0]})));
 assign mul_22_25_n_666 = ~((mul_22_25_n_316 | mul_22_25_n_26) & (mul_22_25_n_590 | mul_22_25_n_292));
 assign mul_22_25_n_665 = ~((mul_22_25_n_277 | mul_22_25_n_26) & (mul_22_25_n_590 | mul_22_25_n_251));
 assign mul_22_25_n_688 = ~(mul_22_25_n_591 & (mul_22_25_n_590 | mul_22_25_n_568));
 assign mul_22_25_n_687 = ~((mul_22_25_n_382 & {in2[0]}) | (mul_22_25_n_589 & mul_22_25_n_70));
 assign mul_22_25_n_686 = ~(mul_22_25_n_591 & (mul_22_25_n_590 | mul_22_25_n_561));
 assign mul_22_25_n_685 = ~((mul_22_25_n_425 & {in2[0]}) | (mul_22_25_n_589 & mul_22_25_n_317));
 assign mul_22_25_n_656 = ~((mul_22_25_n_251 | mul_22_25_n_26) & (mul_22_25_n_590 | mul_22_25_n_234));
 assign mul_22_25_n_655 = ~((mul_22_25_n_249 | mul_22_25_n_26) & (mul_22_25_n_590 | mul_22_25_n_293));
 assign mul_22_25_n_654 = ~((mul_22_25_n_489 | mul_22_25_n_26) & (mul_22_25_n_590 | mul_22_25_n_504));
 assign mul_22_25_n_653 = ~((mul_22_25_n_479 | mul_22_25_n_26) & (mul_22_25_n_590 | mul_22_25_n_437));
 assign mul_22_25_n_652 = ~((mul_22_25_n_561 | mul_22_25_n_26) & (mul_22_25_n_590 | mul_22_25_n_550));
 assign mul_22_25_n_651 = ~((mul_22_25_n_527 | mul_22_25_n_26) & (mul_22_25_n_590 | mul_22_25_n_489));
 assign mul_22_25_n_650 = ~((mul_22_25_n_376 | mul_22_25_n_26) & (mul_22_25_n_590 | mul_22_25_n_277));
 assign mul_22_25_n_649 = ~((mul_22_25_n_236 | mul_22_25_n_26) & (mul_22_25_n_590 | mul_22_25_n_376));
 assign mul_22_25_n_648 = ~((mul_22_25_n_304 | mul_22_25_n_26) & (mul_22_25_n_590 | mul_22_25_n_236));
 assign mul_22_25_n_647 = ((mul_22_25_n_442 & {in2[0]}) | (mul_22_25_n_589 & mul_22_25_n_425));
 assign mul_22_25_n_646 = ~((mul_22_25_n_547 | mul_22_25_n_26) & (mul_22_25_n_590 | mul_22_25_n_526));
 assign mul_22_25_n_645 = ~((mul_22_25_n_437 | mul_22_25_n_26) & (mul_22_25_n_590 | mul_22_25_n_441));
 assign mul_22_25_n_644 = ~((mul_22_25_n_93 | mul_22_25_n_26) & (mul_22_25_n_590 | mul_22_25_n_244));
 assign mul_22_25_n_643 = ~((mul_22_25_n_407 | mul_22_25_n_26) & (mul_22_25_n_590 | mul_22_25_n_260));
 assign mul_22_25_n_642 = ~((mul_22_25_n_299 | mul_22_25_n_26) & (mul_22_25_n_590 | mul_22_25_n_256));
 assign mul_22_25_n_641 = ~((mul_22_25_n_468 | mul_22_25_n_26) & (mul_22_25_n_590 | mul_22_25_n_479));
 assign mul_22_25_n_664 = ~((mul_22_25_n_232 & {in2[0]}) | (mul_22_25_n_589 & mul_22_25_n_382));
 assign mul_22_25_n_663 = ~((~mul_22_25_n_292 & ~mul_22_25_n_26) | (mul_22_25_n_589 & mul_22_25_n_298));
 assign mul_22_25_n_662 = ~((mul_22_25_n_294 & {in2[0]}) | (mul_22_25_n_589 & mul_22_25_n_92));
 assign mul_22_25_n_661 = ~((mul_22_25_n_261 & {in2[0]}) | (mul_22_25_n_589 & mul_22_25_n_305));
 assign mul_22_25_n_660 = ~((mul_22_25_n_243 & {in2[0]}) | (mul_22_25_n_589 & mul_22_25_n_232));
 assign mul_22_25_n_659 = ~((mul_22_25_n_255 & {in2[0]}) | (mul_22_25_n_589 & mul_22_25_n_408));
 assign mul_22_25_n_658 = ~((mul_22_25_n_549 & {in2[0]}) | (mul_22_25_n_589 & mul_22_25_n_546));
 assign mul_22_25_n_657 = ~((mul_22_25_n_235 & {in2[0]}) | (mul_22_25_n_589 & mul_22_25_n_250));
 assign mul_22_25_n_639 = ~mul_22_25_n_3;
 assign mul_22_25_n_638 = ~mul_22_25_n_5;
 assign mul_22_25_n_636 = ~(mul_22_25_n_362 | mul_22_25_n_23);
 assign mul_22_25_n_635 = ~(mul_22_25_n_354 | mul_22_25_n_23);
 assign mul_22_25_n_634 = ~(mul_22_25_n_349 | mul_22_25_n_23);
 assign mul_22_25_n_633 = ~(mul_22_25_n_363 | mul_22_25_n_23);
 assign mul_22_25_n_632 = ~(mul_22_25_n_357 | mul_22_25_n_23);
 assign mul_22_25_n_631 = ~(mul_22_25_n_361 | mul_22_25_n_23);
 assign mul_22_25_n_630 = ~(mul_22_25_n_353 | mul_22_25_n_23);
 assign mul_22_25_n_629 = ~(mul_22_25_n_358 | mul_22_25_n_23);
 assign mul_22_25_n_628 = ~(mul_22_25_n_352 | mul_22_25_n_23);
 assign mul_22_25_n_627 = ~(mul_22_25_n_350 | mul_22_25_n_23);
 assign mul_22_25_n_626 = ~(mul_22_25_n_356 | mul_22_25_n_23);
 assign mul_22_25_n_625 = ~(mul_22_25_n_359 | mul_22_25_n_23);
 assign mul_22_25_n_624 = ~(mul_22_25_n_355 | mul_22_25_n_23);
 assign mul_22_25_n_623 = ~(mul_22_25_n_360 | mul_22_25_n_23);
 assign mul_22_25_n_640 = (mul_22_25_n_593 & mul_22_25_n_560);
 assign mul_22_25_n_637 = ~(mul_22_25_n_594 & {in1[0]});
 assign mul_22_25_n_622 = ~mul_22_25_n_6;
 assign mul_22_25_n_621 = ~mul_22_25_n_7;
 assign mul_22_25_n_620 = ~mul_22_25_n_4;
 assign mul_22_25_n_611 = ~mul_22_25_n_612;
 assign mul_22_25_n_609 = ~mul_22_25_n_610;
 assign mul_22_25_n_607 = ~mul_22_25_n_608;
 assign mul_22_25_n_605 = ~mul_22_25_n_606;
 assign mul_22_25_n_603 = ~mul_22_25_n_604;
 assign mul_22_25_n_601 = ~mul_22_25_n_602;
 assign mul_22_25_n_599 = ~mul_22_25_n_600;
 assign mul_22_25_n_597 = ~mul_22_25_n_598;
 assign mul_22_25_n_595 = ~mul_22_25_n_596;
 assign mul_22_25_n_619 = (mul_22_25_n_594 & mul_22_25_n_559);
 assign mul_22_25_n_618 = ~(mul_22_25_n_363 & mul_22_25_n_334);
 assign mul_22_25_n_617 = ~(mul_22_25_n_362 & mul_22_25_n_335);
 assign mul_22_25_n_616 = ~(mul_22_25_n_361 & mul_22_25_n_336);
 assign mul_22_25_n_615 = ~(mul_22_25_n_360 & mul_22_25_n_337);
 assign mul_22_25_n_614 = ~(mul_22_25_n_359 & mul_22_25_n_338);
 assign mul_22_25_n_613 = ~(mul_22_25_n_358 & mul_22_25_n_339);
 assign mul_22_25_n_612 = ~(mul_22_25_n_354 & mul_22_25_n_345);
 assign mul_22_25_n_610 = ~(mul_22_25_n_353 & mul_22_25_n_346);
 assign mul_22_25_n_608 = ~(mul_22_25_n_357 & mul_22_25_n_348);
 assign mul_22_25_n_606 = ~(mul_22_25_n_350 & mul_22_25_n_344);
 assign mul_22_25_n_604 = ~(mul_22_25_n_352 & mul_22_25_n_347);
 assign mul_22_25_n_602 = ~(mul_22_25_n_349 & mul_22_25_n_343);
 assign mul_22_25_n_600 = ~(mul_22_25_n_356 & mul_22_25_n_340);
 assign mul_22_25_n_598 = ~(mul_22_25_n_355 & mul_22_25_n_341);
 assign mul_22_25_n_596 = ~(mul_22_25_n_351 & mul_22_25_n_342);
 assign mul_22_25_n_594 = ~mul_22_25_n_351;
 assign mul_22_25_n_593 = ~mul_22_25_n_349;
 assign mul_22_25_n_592 = ~mul_22_25_n_354;
 assign mul_22_25_n_591 = ~({in2[0]} & ~mul_22_25_n_568);
 assign mul_22_25_n_589 = ~mul_22_25_n_590;
 assign mul_22_25_n_590 = ~({in2[1]} & mul_22_25_n_26);
 assign mul_22_25_n_557 = ~mul_22_25_n_556;
 assign mul_22_25_n_552 = ~mul_22_25_n_551;
 assign mul_22_25_n_550 = ~mul_22_25_n_549;
 assign mul_22_25_n_547 = ~mul_22_25_n_546;
 assign mul_22_25_n_538 = ~mul_22_25_n_537;
 assign mul_22_25_n_472 = ~mul_22_25_n_471;
 assign mul_22_25_n_450 = ~mul_22_25_n_449;
 assign mul_22_25_n_442 = ~mul_22_25_n_441;
 assign mul_22_25_n_408 = ~mul_22_25_n_407;
 assign mul_22_25_n_348 = ~((mul_22_25_n_18 & ~{in2[10]}) | ({in2[11]} & {in2[10]}));
 assign mul_22_25_n_347 = ~((mul_22_25_n_43 & ~{in2[4]}) | ({in2[5]} & {in2[4]}));
 assign mul_22_25_n_346 = ~((mul_22_25_n_40 & ~{in2[16]}) | ({in2[17]} & {in2[16]}));
 assign mul_22_25_n_345 = ~((mul_22_25_n_41 & ~{in2[18]}) | ({in2[19]} & {in2[18]}));
 assign mul_22_25_n_344 = ~((mul_22_25_n_19 & ~{in2[14]}) | ({in2[15]} & {in2[14]}));
 assign mul_22_25_n_343 = ~((mul_22_25_n_21 & ~{in2[12]}) | ({in2[13]} & {in2[12]}));
 assign mul_22_25_n_342 = ~((mul_22_25_n_42 & ~{in2[2]}) | ({in2[3]} & {in2[2]}));
 assign mul_22_25_n_341 = ~((mul_22_25_n_20 & ~{in2[6]}) | ({in2[7]} & {in2[6]}));
 assign mul_22_25_n_340 = ~((mul_22_25_n_17 & ~{in2[8]}) | ({in2[9]} & {in2[8]}));
 assign mul_22_25_n_339 = ~((mul_22_25_n_22 & ~{in2[20]}) | ({in2[21]} & {in2[20]}));
 assign mul_22_25_n_338 = ~((mul_22_25_n_45 & ~{in2[22]}) | ({in2[23]} & {in2[22]}));
 assign mul_22_25_n_337 = ~((mul_22_25_n_24 & ~{in2[24]}) | ({in2[25]} & {in2[24]}));
 assign mul_22_25_n_336 = ~((mul_22_25_n_25 & ~{in2[26]}) | ({in2[27]} & {in2[26]}));
 assign mul_22_25_n_335 = ~((mul_22_25_n_46 & ~{in2[28]}) | ({in2[29]} & {in2[28]}));
 assign mul_22_25_n_334 = ~((mul_22_25_n_47 & ~{in2[30]}) | ({in2[31]} & {in2[30]}));
 assign mul_22_25_n_333 = ~(({in1[31]} | mul_22_25_n_41) & ({in2[19]} | mul_22_25_n_38));
 assign mul_22_25_n_332 = ~((mul_22_25_n_65 & {in2[21]}) | (mul_22_25_n_22 & {in1[29]}));
 assign mul_22_25_n_331 = ~((mul_22_25_n_63 & {in2[23]}) | (mul_22_25_n_45 & {in1[27]}));
 assign mul_22_25_n_330 = ~((mul_22_25_n_62 & {in2[25]}) | (mul_22_25_n_24 & {in1[25]}));
 assign mul_22_25_n_329 = ~((mul_22_25_n_34 & {in2[27]}) | (mul_22_25_n_25 & {in1[23]}));
 assign mul_22_25_n_588 = ~((mul_22_25_n_61 & {in2[19]}) | (mul_22_25_n_41 & {in1[14]}));
 assign mul_22_25_n_587 = ~((mul_22_25_n_60 & {in2[15]}) | (mul_22_25_n_19 & {in1[18]}));
 assign mul_22_25_n_586 = ~((mul_22_25_n_49 & {in2[17]}) | (mul_22_25_n_40 & {in1[12]}));
 assign mul_22_25_n_585 = ~((mul_22_25_n_54 & {in2[3]}) | (mul_22_25_n_42 & {in1[1]}));
 assign mul_22_25_n_584 = ~((mul_22_25_n_58 & {in2[7]}) | (mul_22_25_n_20 & {in1[8]}));
 assign mul_22_25_n_583 = ~((mul_22_25_n_61 & {in2[11]}) | (mul_22_25_n_18 & {in1[14]}));
 assign mul_22_25_n_582 = ~((mul_22_25_n_54 & {in2[5]}) | (mul_22_25_n_43 & {in1[1]}));
 assign mul_22_25_n_581 = ~((mul_22_25_n_59 & {in2[9]}) | (mul_22_25_n_17 & {in1[2]}));
 assign mul_22_25_n_580 = ~((mul_22_25_n_58 & {in2[13]}) | (mul_22_25_n_21 & {in1[8]}));
 assign mul_22_25_n_579 = ~((mul_22_25_n_55 & {in2[17]}) | (mul_22_25_n_40 & {in1[15]}));
 assign mul_22_25_n_578 = ~((mul_22_25_n_56 & {in2[11]}) | (mul_22_25_n_18 & {in1[13]}));
 assign mul_22_25_n_577 = ~(({in1[30]} | mul_22_25_n_41) & ({in2[19]} | mul_22_25_n_39));
 assign mul_22_25_n_576 = ~(({in1[30]} | mul_22_25_n_42) & ({in2[3]} | mul_22_25_n_39));
 assign mul_22_25_n_575 = ~(({in1[31]} | mul_22_25_n_40) & ({in2[17]} | mul_22_25_n_38));
 assign mul_22_25_n_574 = ~((mul_22_25_n_39 & {in2[9]}) | (mul_22_25_n_17 & {in1[30]}));
 assign mul_22_25_n_573 = ~((mul_22_25_n_39 & {in2[13]}) | (mul_22_25_n_21 & {in1[30]}));
 assign mul_22_25_n_572 = ~(({in1[31]} | mul_22_25_n_43) & ({in2[5]} | mul_22_25_n_38));
 assign mul_22_25_n_571 = ~((mul_22_25_n_50 & {in2[13]}) | (mul_22_25_n_21 & {in1[17]}));
 assign mul_22_25_n_570 = ~(({in1[31]} | mul_22_25_n_17) & ({in2[9]} | mul_22_25_n_38));
 assign mul_22_25_n_569 = ~((mul_22_25_n_39 & {in2[11]}) | (mul_22_25_n_18 & {in1[30]}));
 assign mul_22_25_n_568 = ~((mul_22_25_n_38 & {in2[1]}) | (mul_22_25_n_44 & {in1[31]}));
 assign mul_22_25_n_567 = ~(({in1[31]} | mul_22_25_n_19) & ({in2[15]} | mul_22_25_n_38));
 assign mul_22_25_n_566 = ~(({in1[31]} | mul_22_25_n_20) & ({in2[7]} | mul_22_25_n_38));
 assign mul_22_25_n_565 = ~(({in1[31]} | mul_22_25_n_18) & ({in2[11]} | mul_22_25_n_38));
 assign mul_22_25_n_564 = ~((mul_22_25_n_39 & {in2[7]}) | (mul_22_25_n_20 & {in1[30]}));
 assign mul_22_25_n_563 = ~((mul_22_25_n_39 & {in2[17]}) | (mul_22_25_n_40 & {in1[30]}));
 assign mul_22_25_n_562 = ~((mul_22_25_n_39 & {in2[15]}) | (mul_22_25_n_19 & {in1[30]}));
 assign mul_22_25_n_561 = ~((mul_22_25_n_39 & {in2[1]}) | (mul_22_25_n_44 & {in1[30]}));
 assign mul_22_25_n_560 = ~(({in1[31]} | mul_22_25_n_21) & ({in2[13]} | mul_22_25_n_38));
 assign mul_22_25_n_559 = ~(({in1[31]} | mul_22_25_n_42) & ({in2[3]} | mul_22_25_n_38));
 assign mul_22_25_n_558 = ~((mul_22_25_n_39 & {in2[5]}) | (mul_22_25_n_43 & {in1[30]}));
 assign mul_22_25_n_556 = ~((mul_22_25_n_64 & {in2[13]}) | (mul_22_25_n_21 & {in1[28]}));
 assign mul_22_25_n_555 = ~((mul_22_25_n_65 & {in2[5]}) | (mul_22_25_n_43 & {in1[29]}));
 assign mul_22_25_n_554 = ~((mul_22_25_n_64 & {in2[9]}) | (mul_22_25_n_17 & {in1[28]}));
 assign mul_22_25_n_553 = ~((mul_22_25_n_65 & {in2[17]}) | (mul_22_25_n_40 & {in1[29]}));
 assign mul_22_25_n_551 = ~((mul_22_25_n_65 & {in2[13]}) | (mul_22_25_n_21 & {in1[29]}));
 assign mul_22_25_n_549 = ~(({in1[29]} | mul_22_25_n_44) & ({in2[1]} | mul_22_25_n_65));
 assign mul_22_25_n_548 = ~((mul_22_25_n_64 & {in2[19]}) | (mul_22_25_n_41 & {in1[28]}));
 assign mul_22_25_n_546 = ~(({in1[28]} | mul_22_25_n_44) & ({in2[1]} | mul_22_25_n_64));
 assign mul_22_25_n_545 = ~((mul_22_25_n_65 & {in2[3]}) | (mul_22_25_n_42 & {in1[29]}));
 assign mul_22_25_n_544 = ~((mul_22_25_n_64 & {in2[11]}) | (mul_22_25_n_18 & {in1[28]}));
 assign mul_22_25_n_543 = ~((mul_22_25_n_64 & {in2[5]}) | (mul_22_25_n_43 & {in1[28]}));
 assign mul_22_25_n_542 = ~((mul_22_25_n_64 & {in2[3]}) | (mul_22_25_n_42 & {in1[28]}));
 assign mul_22_25_n_541 = ~((mul_22_25_n_64 & {in2[15]}) | (mul_22_25_n_19 & {in1[28]}));
 assign mul_22_25_n_540 = ~((mul_22_25_n_65 & {in2[15]}) | (mul_22_25_n_19 & {in1[29]}));
 assign mul_22_25_n_539 = ~((mul_22_25_n_65 & {in2[7]}) | (mul_22_25_n_20 & {in1[29]}));
 assign mul_22_25_n_537 = ~((mul_22_25_n_65 & {in2[19]}) | (mul_22_25_n_41 & {in1[29]}));
 assign mul_22_25_n_536 = ~((mul_22_25_n_65 & {in2[9]}) | (mul_22_25_n_17 & {in1[29]}));
 assign mul_22_25_n_535 = ~((mul_22_25_n_65 & {in2[11]}) | (mul_22_25_n_18 & {in1[29]}));
 assign mul_22_25_n_534 = ~((mul_22_25_n_64 & {in2[17]}) | (mul_22_25_n_40 & {in1[28]}));
 assign mul_22_25_n_533 = ~((mul_22_25_n_64 & {in2[7]}) | (mul_22_25_n_20 & {in1[28]}));
 assign mul_22_25_n_532 = ~((mul_22_25_n_60 & {in2[3]}) | (mul_22_25_n_42 & {in1[18]}));
 assign mul_22_25_n_531 = ~((mul_22_25_n_64 & {in2[21]}) | (mul_22_25_n_22 & {in1[28]}));
 assign mul_22_25_n_530 = ~((mul_22_25_n_37 & {in2[17]}) | (mul_22_25_n_40 & {in1[26]}));
 assign mul_22_25_n_529 = ~((mul_22_25_n_63 & {in2[13]}) | (mul_22_25_n_21 & {in1[27]}));
 assign mul_22_25_n_528 = ~((mul_22_25_n_37 & {in2[3]}) | (mul_22_25_n_42 & {in1[26]}));
 assign mul_22_25_n_527 = ~((mul_22_25_n_37 & {in2[1]}) | (mul_22_25_n_44 & {in1[26]}));
 assign mul_22_25_n_526 = ~((mul_22_25_n_63 & {in2[1]}) | (mul_22_25_n_44 & {in1[27]}));
 assign mul_22_25_n_525 = ~((mul_22_25_n_37 & {in2[7]}) | (mul_22_25_n_20 & {in1[26]}));
 assign mul_22_25_n_524 = ~((mul_22_25_n_63 & {in2[7]}) | (mul_22_25_n_20 & {in1[27]}));
 assign mul_22_25_n_523 = ~((mul_22_25_n_63 & {in2[15]}) | (mul_22_25_n_19 & {in1[27]}));
 assign mul_22_25_n_522 = ~((mul_22_25_n_63 & {in2[19]}) | (mul_22_25_n_41 & {in1[27]}));
 assign mul_22_25_n_521 = ~((mul_22_25_n_37 & {in2[5]}) | (mul_22_25_n_43 & {in1[26]}));
 assign mul_22_25_n_520 = ~((mul_22_25_n_37 & {in2[19]}) | (mul_22_25_n_41 & {in1[26]}));
 assign mul_22_25_n_519 = ~((mul_22_25_n_37 & {in2[9]}) | (mul_22_25_n_17 & {in1[26]}));
 assign mul_22_25_n_518 = ~((mul_22_25_n_37 & {in2[15]}) | (mul_22_25_n_19 & {in1[26]}));
 assign mul_22_25_n_517 = ~((mul_22_25_n_63 & {in2[17]}) | (mul_22_25_n_40 & {in1[27]}));
 assign mul_22_25_n_516 = ~((mul_22_25_n_63 & {in2[3]}) | (mul_22_25_n_42 & {in1[27]}));
 assign mul_22_25_n_515 = ~((mul_22_25_n_63 & {in2[9]}) | (mul_22_25_n_17 & {in1[27]}));
 assign mul_22_25_n_514 = ~((mul_22_25_n_63 & {in2[11]}) | (mul_22_25_n_18 & {in1[27]}));
 assign mul_22_25_n_513 = ~((mul_22_25_n_37 & {in2[13]}) | (mul_22_25_n_21 & {in1[26]}));
 assign mul_22_25_n_512 = ~((mul_22_25_n_63 & {in2[5]}) | (mul_22_25_n_43 & {in1[27]}));
 assign mul_22_25_n_511 = ~((mul_22_25_n_37 & {in2[11]}) | (mul_22_25_n_18 & {in1[26]}));
 assign mul_22_25_n_510 = ~((mul_22_25_n_37 & {in2[21]}) | (mul_22_25_n_22 & {in1[26]}));
 assign mul_22_25_n_509 = ~((mul_22_25_n_63 & {in2[21]}) | (mul_22_25_n_22 & {in1[27]}));
 assign mul_22_25_n_508 = ~({in2[1]} & ~asc001_0_);
 assign mul_22_25_n_507 = ~((mul_22_25_n_37 & {in2[23]}) | (mul_22_25_n_45 & {in1[26]}));
 assign mul_22_25_n_506 = ~((mul_22_25_n_36 & {in2[11]}) | (mul_22_25_n_18 & {in1[24]}));
 assign mul_22_25_n_505 = ~((mul_22_25_n_62 & {in2[11]}) | (mul_22_25_n_18 & {in1[25]}));
 assign mul_22_25_n_504 = ~((mul_22_25_n_36 & {in2[1]}) | (mul_22_25_n_44 & {in1[24]}));
 assign mul_22_25_n_503 = ~((mul_22_25_n_36 & {in2[7]}) | (mul_22_25_n_20 & {in1[24]}));
 assign mul_22_25_n_502 = ~((mul_22_25_n_62 & {in2[5]}) | (mul_22_25_n_43 & {in1[25]}));
 assign mul_22_25_n_501 = ~((mul_22_25_n_62 & {in2[13]}) | (mul_22_25_n_21 & {in1[25]}));
 assign mul_22_25_n_500 = ~((mul_22_25_n_36 & {in2[13]}) | (mul_22_25_n_21 & {in1[24]}));
 assign mul_22_25_n_499 = ~((mul_22_25_n_36 & {in2[19]}) | (mul_22_25_n_41 & {in1[24]}));
 assign mul_22_25_n_498 = ~((mul_22_25_n_36 & {in2[3]}) | (mul_22_25_n_42 & {in1[24]}));
 assign mul_22_25_n_497 = ~((mul_22_25_n_36 & {in2[17]}) | (mul_22_25_n_40 & {in1[24]}));
 assign mul_22_25_n_496 = ~((mul_22_25_n_62 & {in2[7]}) | (mul_22_25_n_20 & {in1[25]}));
 assign mul_22_25_n_495 = ~((mul_22_25_n_62 & {in2[9]}) | (mul_22_25_n_17 & {in1[25]}));
 assign mul_22_25_n_494 = ~((mul_22_25_n_62 & {in2[19]}) | (mul_22_25_n_41 & {in1[25]}));
 assign mul_22_25_n_493 = ~((mul_22_25_n_36 & {in2[9]}) | (mul_22_25_n_17 & {in1[24]}));
 assign mul_22_25_n_492 = ~((mul_22_25_n_36 & {in2[15]}) | (mul_22_25_n_19 & {in1[24]}));
 assign mul_22_25_n_491 = ~((mul_22_25_n_62 & {in2[17]}) | (mul_22_25_n_40 & {in1[25]}));
 assign mul_22_25_n_490 = ~((mul_22_25_n_62 & {in2[3]}) | (mul_22_25_n_42 & {in1[25]}));
 assign mul_22_25_n_489 = ~((mul_22_25_n_62 & {in2[1]}) | (mul_22_25_n_44 & {in1[25]}));
 assign mul_22_25_n_488 = ~((mul_22_25_n_36 & {in2[5]}) | (mul_22_25_n_43 & {in1[24]}));
 assign mul_22_25_n_487 = ~((mul_22_25_n_62 & {in2[15]}) | (mul_22_25_n_19 & {in1[25]}));
 assign mul_22_25_n_486 = ~((mul_22_25_n_36 & {in2[21]}) | (mul_22_25_n_22 & {in1[24]}));
 assign mul_22_25_n_485 = ~((mul_22_25_n_62 & {in2[21]}) | (mul_22_25_n_22 & {in1[25]}));
 assign mul_22_25_n_484 = ~((mul_22_25_n_36 & {in2[23]}) | (mul_22_25_n_45 & {in1[24]}));
 assign mul_22_25_n_483 = ~((mul_22_25_n_62 & {in2[23]}) | (mul_22_25_n_45 & {in1[25]}));
 assign mul_22_25_n_482 = ~((mul_22_25_n_35 & {in2[11]}) | (mul_22_25_n_18 & {in1[22]}));
 assign mul_22_25_n_481 = ~((mul_22_25_n_34 & {in2[7]}) | (mul_22_25_n_20 & {in1[23]}));
 assign mul_22_25_n_480 = ~((mul_22_25_n_35 & {in2[7]}) | (mul_22_25_n_20 & {in1[22]}));
 assign mul_22_25_n_479 = ~((mul_22_25_n_35 & {in2[1]}) | (mul_22_25_n_44 & {in1[22]}));
 assign mul_22_25_n_478 = ~((mul_22_25_n_35 & {in2[15]}) | (mul_22_25_n_19 & {in1[22]}));
 assign mul_22_25_n_477 = ~((mul_22_25_n_34 & {in2[9]}) | (mul_22_25_n_17 & {in1[23]}));
 assign mul_22_25_n_476 = ~((mul_22_25_n_35 & {in2[17]}) | (mul_22_25_n_40 & {in1[22]}));
 assign mul_22_25_n_475 = ~((mul_22_25_n_34 & {in2[11]}) | (mul_22_25_n_18 & {in1[23]}));
 assign mul_22_25_n_474 = ~((mul_22_25_n_35 & {in2[19]}) | (mul_22_25_n_41 & {in1[22]}));
 assign mul_22_25_n_473 = ~((mul_22_25_n_34 & {in2[13]}) | (mul_22_25_n_21 & {in1[23]}));
 assign mul_22_25_n_471 = ~((mul_22_25_n_34 & {in2[3]}) | (mul_22_25_n_42 & {in1[23]}));
 assign mul_22_25_n_470 = ~(({in1[22]} | mul_22_25_n_42) & ({in2[3]} | mul_22_25_n_35));
 assign mul_22_25_n_469 = ~((mul_22_25_n_35 & {in2[5]}) | (mul_22_25_n_43 & {in1[22]}));
 assign mul_22_25_n_468 = ~((mul_22_25_n_34 & {in2[1]}) | (mul_22_25_n_44 & {in1[23]}));
 assign mul_22_25_n_467 = ~((mul_22_25_n_34 & {in2[15]}) | (mul_22_25_n_19 & {in1[23]}));
 assign mul_22_25_n_466 = ~((mul_22_25_n_35 & {in2[9]}) | (mul_22_25_n_17 & {in1[22]}));
 assign mul_22_25_n_465 = ~((mul_22_25_n_34 & {in2[19]}) | (mul_22_25_n_41 & {in1[23]}));
 assign mul_22_25_n_464 = ~((mul_22_25_n_34 & {in2[17]}) | (mul_22_25_n_40 & {in1[23]}));
 assign mul_22_25_n_463 = ~((mul_22_25_n_35 & {in2[13]}) | (mul_22_25_n_21 & {in1[22]}));
 assign mul_22_25_n_462 = ~((mul_22_25_n_34 & {in2[5]}) | (mul_22_25_n_43 & {in1[23]}));
 assign mul_22_25_n_461 = ~((mul_22_25_n_36 & {in2[25]}) | (mul_22_25_n_24 & {in1[24]}));
 assign mul_22_25_n_460 = ~((mul_22_25_n_55 & {in2[7]}) | (mul_22_25_n_20 & {in1[15]}));
 assign mul_22_25_n_459 = ~((mul_22_25_n_34 & {in2[21]}) | (mul_22_25_n_22 & {in1[23]}));
 assign mul_22_25_n_458 = ~((mul_22_25_n_35 & {in2[21]}) | (mul_22_25_n_22 & {in1[22]}));
 assign mul_22_25_n_457 = ~((mul_22_25_n_35 & {in2[23]}) | (mul_22_25_n_45 & {in1[22]}));
 assign mul_22_25_n_456 = ~((mul_22_25_n_34 & {in2[23]}) | (mul_22_25_n_45 & {in1[23]}));
 assign mul_22_25_n_455 = ~((mul_22_25_n_32 & {in2[11]}) | (mul_22_25_n_18 & {in1[21]}));
 assign mul_22_25_n_454 = ~((mul_22_25_n_32 & {in2[7]}) | (mul_22_25_n_20 & {in1[21]}));
 assign mul_22_25_n_453 = ~((mul_22_25_n_33 & {in2[17]}) | (mul_22_25_n_40 & {in1[20]}));
 assign mul_22_25_n_452 = ~((mul_22_25_n_32 & {in2[19]}) | (mul_22_25_n_41 & {in1[21]}));
 assign mul_22_25_n_451 = ~((mul_22_25_n_33 & {in2[19]}) | (mul_22_25_n_41 & {in1[20]}));
 assign mul_22_25_n_449 = ~(({in1[21]} | mul_22_25_n_42) & ({in2[3]} | mul_22_25_n_32));
 assign mul_22_25_n_448 = ~((mul_22_25_n_32 & {in2[17]}) | (mul_22_25_n_40 & {in1[21]}));
 assign mul_22_25_n_447 = ~((mul_22_25_n_32 & {in2[13]}) | (mul_22_25_n_21 & {in1[21]}));
 assign mul_22_25_n_446 = ~((mul_22_25_n_32 & {in2[15]}) | (mul_22_25_n_19 & {in1[21]}));
 assign mul_22_25_n_445 = ~((mul_22_25_n_33 & {in2[13]}) | (mul_22_25_n_21 & {in1[20]}));
 assign mul_22_25_n_444 = ~((mul_22_25_n_33 & {in2[3]}) | (mul_22_25_n_42 & {in1[20]}));
 assign mul_22_25_n_443 = ~((mul_22_25_n_33 & {in2[11]}) | (mul_22_25_n_18 & {in1[20]}));
 assign mul_22_25_n_441 = ~((mul_22_25_n_33 & {in2[1]}) | (mul_22_25_n_44 & {in1[20]}));
 assign mul_22_25_n_440 = ~((mul_22_25_n_33 & {in2[15]}) | (mul_22_25_n_19 & {in1[20]}));
 assign mul_22_25_n_439 = ~((mul_22_25_n_33 & {in2[9]}) | (mul_22_25_n_17 & {in1[20]}));
 assign mul_22_25_n_438 = ~((mul_22_25_n_32 & {in2[9]}) | (mul_22_25_n_17 & {in1[21]}));
 assign mul_22_25_n_437 = ~((mul_22_25_n_32 & {in2[1]}) | (mul_22_25_n_44 & {in1[21]}));
 assign mul_22_25_n_436 = ~((mul_22_25_n_33 & {in2[7]}) | (mul_22_25_n_20 & {in1[20]}));
 assign mul_22_25_n_435 = ~((mul_22_25_n_33 & {in2[5]}) | (mul_22_25_n_43 & {in1[20]}));
 assign mul_22_25_n_434 = ~((mul_22_25_n_32 & {in2[5]}) | (mul_22_25_n_43 & {in1[21]}));
 assign mul_22_25_n_433 = ~((mul_22_25_n_35 & {in2[25]}) | (mul_22_25_n_24 & {in1[22]}));
 assign mul_22_25_n_432 = ~((mul_22_25_n_34 & {in2[25]}) | (mul_22_25_n_24 & {in1[23]}));
 assign mul_22_25_n_431 = ~((mul_22_25_n_33 & {in2[21]}) | (mul_22_25_n_22 & {in1[20]}));
 assign mul_22_25_n_430 = ~((mul_22_25_n_32 & {in2[21]}) | (mul_22_25_n_22 & {in1[21]}));
 assign mul_22_25_n_429 = ~((mul_22_25_n_35 & {in2[27]}) | (mul_22_25_n_25 & {in1[22]}));
 assign mul_22_25_n_428 = ~(({in1[6]} | mul_22_25_n_42) & ({in2[3]} | mul_22_25_n_52));
 assign mul_22_25_n_427 = ~((mul_22_25_n_33 & {in2[23]}) | (mul_22_25_n_45 & {in1[20]}));
 assign mul_22_25_n_426 = ~((mul_22_25_n_32 & {in2[23]}) | (mul_22_25_n_45 & {in1[21]}));
 assign mul_22_25_n_425 = ~(({in1[19]} | mul_22_25_n_44) & ({in2[1]} | mul_22_25_n_48));
 assign mul_22_25_n_424 = ~((mul_22_25_n_52 & {in2[15]}) | (mul_22_25_n_19 & {in1[6]}));
 assign mul_22_25_n_423 = ~((mul_22_25_n_52 & {in2[5]}) | (mul_22_25_n_43 & {in1[6]}));
 assign mul_22_25_n_422 = ~((mul_22_25_n_28 & {in2[11]}) | (mul_22_25_n_18 & {in1[3]}));
 assign mul_22_25_n_421 = ~((mul_22_25_n_30 & {in2[19]}) | (mul_22_25_n_41 & {in1[4]}));
 assign mul_22_25_n_420 = ~((mul_22_25_n_60 & {in2[7]}) | (mul_22_25_n_20 & {in1[18]}));
 assign mul_22_25_n_419 = ~((mul_22_25_n_57 & {in2[19]}) | (mul_22_25_n_41 & {in1[5]}));
 assign mul_22_25_n_418 = ~((mul_22_25_n_56 & {in2[13]}) | (mul_22_25_n_21 & {in1[13]}));
 assign mul_22_25_n_417 = ~((mul_22_25_n_61 & {in2[13]}) | (mul_22_25_n_21 & {in1[14]}));
 assign mul_22_25_n_416 = ~((mul_22_25_n_51 & {in2[9]}) | (mul_22_25_n_17 & {in1[16]}));
 assign mul_22_25_n_415 = ~((mul_22_25_n_51 & {in2[13]}) | (mul_22_25_n_21 & {in1[16]}));
 assign mul_22_25_n_414 = ~((mul_22_25_n_59 & {in2[5]}) | (mul_22_25_n_43 & {in1[2]}));
 assign mul_22_25_n_413 = ~((mul_22_25_n_30 & {in2[7]}) | (mul_22_25_n_20 & {in1[4]}));
 assign mul_22_25_n_412 = ~((mul_22_25_n_27 & {in2[17]}) | (mul_22_25_n_40 & {in1[11]}));
 assign mul_22_25_n_411 = ~((mul_22_25_n_54 & {in2[17]}) | (mul_22_25_n_40 & {in1[1]}));
 assign mul_22_25_n_410 = ~((mul_22_25_n_56 & {in2[15]}) | (mul_22_25_n_19 & {in1[13]}));
 assign mul_22_25_n_409 = ~((mul_22_25_n_27 & {in2[9]}) | (mul_22_25_n_17 & {in1[11]}));
 assign mul_22_25_n_407 = ~((mul_22_25_n_61 & {in2[1]}) | (mul_22_25_n_44 & {in1[14]}));
 assign mul_22_25_n_406 = ~(({in1[7]} | mul_22_25_n_42) & ({in2[3]} | mul_22_25_n_31));
 assign mul_22_25_n_405 = ~((mul_22_25_n_49 & {in2[11]}) | (mul_22_25_n_18 & {in1[12]}));
 assign mul_22_25_n_404 = ~((mul_22_25_n_48 & {in2[11]}) | (mul_22_25_n_18 & {in1[19]}));
 assign mul_22_25_n_403 = ~((mul_22_25_n_48 & {in2[3]}) | (mul_22_25_n_42 & {in1[19]}));
 assign mul_22_25_n_402 = ~((mul_22_25_n_61 & {in2[9]}) | (mul_22_25_n_17 & {in1[14]}));
 assign mul_22_25_n_401 = ~((mul_22_25_n_52 & {in2[7]}) | (mul_22_25_n_20 & {in1[6]}));
 assign mul_22_25_n_400 = ~((mul_22_25_n_57 & {in2[13]}) | (mul_22_25_n_21 & {in1[5]}));
 assign mul_22_25_n_399 = ~((mul_22_25_n_30 & {in2[17]}) | (mul_22_25_n_40 & {in1[4]}));
 assign mul_22_25_n_398 = ~((mul_22_25_n_61 & {in2[5]}) | (mul_22_25_n_43 & {in1[14]}));
 assign mul_22_25_n_397 = ~((mul_22_25_n_58 & {in2[9]}) | (mul_22_25_n_17 & {in1[8]}));
 assign mul_22_25_n_396 = ~((mul_22_25_n_27 & {in2[13]}) | (mul_22_25_n_21 & {in1[11]}));
 assign mul_22_25_n_395 = ~((mul_22_25_n_57 & {in2[17]}) | (mul_22_25_n_40 & {in1[5]}));
 assign mul_22_25_n_394 = ~((mul_22_25_n_58 & {in2[17]}) | (mul_22_25_n_40 & {in1[8]}));
 assign mul_22_25_n_393 = ~((mul_22_25_n_55 & {in2[13]}) | (mul_22_25_n_21 & {in1[15]}));
 assign mul_22_25_n_392 = ~((mul_22_25_n_28 & {in2[5]}) | (mul_22_25_n_43 & {in1[3]}));
 assign mul_22_25_n_391 = ~((mul_22_25_n_28 & {in2[3]}) | (mul_22_25_n_42 & {in1[3]}));
 assign mul_22_25_n_390 = ~((mul_22_25_n_48 & {in2[17]}) | (mul_22_25_n_40 & {in1[19]}));
 assign mul_22_25_n_389 = ~((mul_22_25_n_30 & {in2[15]}) | (mul_22_25_n_19 & {in1[4]}));
 assign mul_22_25_n_388 = ~((mul_22_25_n_61 & {in2[17]}) | (mul_22_25_n_40 & {in1[14]}));
 assign mul_22_25_n_387 = ~((mul_22_25_n_31 & {in2[5]}) | (mul_22_25_n_43 & {in1[7]}));
 assign mul_22_25_n_386 = ~((mul_22_25_n_48 & {in2[9]}) | (mul_22_25_n_17 & {in1[19]}));
 assign mul_22_25_n_385 = ~((mul_22_25_n_51 & {in2[17]}) | (mul_22_25_n_40 & {in1[16]}));
 assign mul_22_25_n_384 = ~((mul_22_25_n_58 & {in2[5]}) | (mul_22_25_n_43 & {in1[8]}));
 assign mul_22_25_n_383 = ~((mul_22_25_n_31 & {in2[17]}) | (mul_22_25_n_40 & {in1[7]}));
 assign mul_22_25_n_382 = ~(({in1[1]} | mul_22_25_n_44) & ({in2[1]} | mul_22_25_n_54));
 assign mul_22_25_n_381 = ~((mul_22_25_n_27 & {in2[7]}) | (mul_22_25_n_20 & {in1[11]}));
 assign mul_22_25_n_380 = ~((mul_22_25_n_28 & {in2[15]}) | (mul_22_25_n_19 & {in1[3]}));
 assign mul_22_25_n_379 = ~((mul_22_25_n_55 & {in2[3]}) | (mul_22_25_n_42 & {in1[15]}));
 assign mul_22_25_n_378 = ~((mul_22_25_n_57 & {in2[11]}) | (mul_22_25_n_18 & {in1[5]}));
 assign mul_22_25_n_377 = ~((mul_22_25_n_28 & {in2[17]}) | (mul_22_25_n_40 & {in1[3]}));
 assign mul_22_25_n_376 = ~((mul_22_25_n_53 & {in2[1]}) | (mul_22_25_n_44 & {in1[10]}));
 assign mul_22_25_n_375 = ~((mul_22_25_n_53 & {in2[11]}) | (mul_22_25_n_18 & {in1[10]}));
 assign mul_22_25_n_374 = ~((mul_22_25_n_60 & {in2[13]}) | (mul_22_25_n_21 & {in1[18]}));
 assign mul_22_25_n_373 = ~((mul_22_25_n_60 & {in2[19]}) | (mul_22_25_n_41 & {in1[18]}));
 assign mul_22_25_n_372 = ~((mul_22_25_n_61 & {in2[7]}) | (mul_22_25_n_20 & {in1[14]}));
 assign mul_22_25_n_371 = ~((mul_22_25_n_54 & {in2[9]}) | (mul_22_25_n_17 & {in1[1]}));
 assign mul_22_25_n_370 = ~((mul_22_25_n_51 & {in2[15]}) | (mul_22_25_n_19 & {in1[16]}));
 assign mul_22_25_n_369 = ~((mul_22_25_n_55 & {in2[5]}) | (mul_22_25_n_43 & {in1[15]}));
 assign mul_22_25_n_368 = ~((mul_22_25_n_53 & {in2[3]}) | (mul_22_25_n_42 & {in1[10]}));
 assign mul_22_25_n_367 = ~((mul_22_25_n_53 & {in2[15]}) | (mul_22_25_n_19 & {in1[10]}));
 assign mul_22_25_n_366 = ~((mul_22_25_n_28 & {in2[19]}) | (mul_22_25_n_41 & {in1[3]}));
 assign mul_22_25_n_365 = ~((mul_22_25_n_56 & {in2[3]}) | (mul_22_25_n_42 & {in1[13]}));
 assign mul_22_25_n_364 = ~((mul_22_25_n_31 & {in2[13]}) | (mul_22_25_n_21 & {in1[7]}));
 assign mul_22_25_n_363 = ((mul_22_25_n_46 & ~{in2[30]}) | ({in2[29]} & {in2[30]}));
 assign mul_22_25_n_362 = ((mul_22_25_n_25 & ~{in2[28]}) | ({in2[27]} & {in2[28]}));
 assign mul_22_25_n_361 = ((mul_22_25_n_24 & ~{in2[26]}) | ({in2[25]} & {in2[26]}));
 assign mul_22_25_n_360 = ((mul_22_25_n_45 & ~{in2[24]}) | ({in2[23]} & {in2[24]}));
 assign mul_22_25_n_359 = ((mul_22_25_n_22 & ~{in2[22]}) | ({in2[21]} & {in2[22]}));
 assign mul_22_25_n_358 = ((mul_22_25_n_41 & ~{in2[20]}) | ({in2[19]} & {in2[20]}));
 assign mul_22_25_n_357 = ((mul_22_25_n_17 & ~{in2[10]}) | ({in2[9]} & {in2[10]}));
 assign mul_22_25_n_356 = ((mul_22_25_n_20 & ~{in2[8]}) | ({in2[7]} & {in2[8]}));
 assign mul_22_25_n_355 = ((mul_22_25_n_43 & ~{in2[6]}) | ({in2[5]} & {in2[6]}));
 assign mul_22_25_n_354 = ((mul_22_25_n_40 & ~{in2[18]}) | ({in2[17]} & {in2[18]}));
 assign mul_22_25_n_353 = ((mul_22_25_n_19 & ~{in2[16]}) | ({in2[15]} & {in2[16]}));
 assign mul_22_25_n_352 = ((mul_22_25_n_42 & ~{in2[4]}) | ({in2[3]} & {in2[4]}));
 assign mul_22_25_n_351 = ((mul_22_25_n_44 & ~{in2[2]}) | ({in2[1]} & {in2[2]}));
 assign mul_22_25_n_350 = ((mul_22_25_n_21 & ~{in2[14]}) | ({in2[13]} & {in2[14]}));
 assign mul_22_25_n_349 = ((mul_22_25_n_18 & ~{in2[12]}) | ({in2[11]} & {in2[12]}));
 assign mul_22_25_n_317 = ~mul_22_25_n_316;
 assign mul_22_25_n_305 = ~mul_22_25_n_304;
 assign mul_22_25_n_299 = ~mul_22_25_n_298;
 assign mul_22_25_n_294 = ~mul_22_25_n_293;
 assign mul_22_25_n_261 = ~mul_22_25_n_260;
 assign mul_22_25_n_256 = ~mul_22_25_n_255;
 assign mul_22_25_n_250 = ~mul_22_25_n_249;
 assign mul_22_25_n_244 = ~mul_22_25_n_243;
 assign mul_22_25_n_240 = ~mul_22_25_n_239;
 assign mul_22_25_n_235 = ~mul_22_25_n_234;
 assign mul_22_25_n_93 = ~mul_22_25_n_92;
 assign mul_22_25_n_85 = ~((mul_22_25_n_23 & {in2[17]}) | (mul_22_25_n_40 & {in1[0]}));
 assign mul_22_25_n_84 = ~((mul_22_25_n_32 & {in2[29]}) | (mul_22_25_n_46 & {in1[21]}));
 assign mul_22_25_n_83 = ~((mul_22_25_n_48 & {in2[31]}) | (mul_22_25_n_47 & {in1[19]}));
 assign mul_22_25_n_82 = ~((mul_22_25_n_23 & {in2[31]}) | (mul_22_25_n_47 & {in1[0]}));
 assign mul_22_25_n_81 = ~((mul_22_25_n_23 & {in2[29]}) | (mul_22_25_n_46 & {in1[0]}));
 assign mul_22_25_n_80 = ~((mul_22_25_n_23 & {in2[27]}) | (mul_22_25_n_25 & {in1[0]}));
 assign mul_22_25_n_79 = ~((mul_22_25_n_23 & {in2[9]}) | (mul_22_25_n_17 & {in1[0]}));
 assign mul_22_25_n_78 = ~((mul_22_25_n_23 & {in2[7]}) | (mul_22_25_n_20 & {in1[0]}));
 assign mul_22_25_n_77 = ~((mul_22_25_n_23 & {in2[11]}) | (mul_22_25_n_18 & {in1[0]}));
 assign mul_22_25_n_75 = ~((mul_22_25_n_23 & {in2[19]}) | (mul_22_25_n_41 & {in1[0]}));
 assign mul_22_25_n_74 = ~((mul_22_25_n_23 & {in2[5]}) | (mul_22_25_n_43 & {in1[0]}));
 assign mul_22_25_n_73 = ~((mul_22_25_n_23 & {in2[15]}) | (mul_22_25_n_19 & {in1[0]}));
 assign mul_22_25_n_72 = ~((mul_22_25_n_23 & {in2[3]}) | (mul_22_25_n_42 & {in1[0]}));
 assign mul_22_25_n_71 = ~((mul_22_25_n_23 & {in2[13]}) | (mul_22_25_n_21 & {in1[0]}));
 assign mul_22_25_n_70 = ~(({in1[0]} | mul_22_25_n_44) & ({in2[1]} | mul_22_25_n_23));
 assign mul_22_25_n_69 = ~((mul_22_25_n_23 & {in2[25]}) | (mul_22_25_n_24 & {in1[0]}));
 assign mul_22_25_n_68 = ~((mul_22_25_n_23 & {in2[21]}) | (mul_22_25_n_22 & {in1[0]}));
 assign mul_22_25_n_67 = ~((mul_22_25_n_23 & {in2[23]}) | (mul_22_25_n_45 & {in1[0]}));
 assign mul_22_25_n_328 = ~((mul_22_25_n_60 & {in2[11]}) | (mul_22_25_n_18 & {in1[18]}));
 assign mul_22_25_n_327 = ~((mul_22_25_n_29 & {in2[19]}) | (mul_22_25_n_41 & {in1[9]}));
 assign mul_22_25_n_326 = ~((mul_22_25_n_29 & {in2[13]}) | (mul_22_25_n_21 & {in1[9]}));
 assign mul_22_25_n_325 = ~((mul_22_25_n_59 & {in2[11]}) | (mul_22_25_n_18 & {in1[2]}));
 assign mul_22_25_n_324 = ~((mul_22_25_n_58 & {in2[11]}) | (mul_22_25_n_18 & {in1[8]}));
 assign mul_22_25_n_323 = ~((mul_22_25_n_57 & {in2[7]}) | (mul_22_25_n_20 & {in1[5]}));
 assign mul_22_25_n_322 = ~((mul_22_25_n_58 & {in2[19]}) | (mul_22_25_n_41 & {in1[8]}));
 assign mul_22_25_n_321 = ~((mul_22_25_n_59 & {in2[17]}) | (mul_22_25_n_40 & {in1[2]}));
 assign mul_22_25_n_320 = ~((mul_22_25_n_49 & {in2[15]}) | (mul_22_25_n_19 & {in1[12]}));
 assign mul_22_25_n_319 = ~((mul_22_25_n_53 & {in2[17]}) | (mul_22_25_n_40 & {in1[10]}));
 assign mul_22_25_n_318 = ~((mul_22_25_n_56 & {in2[19]}) | (mul_22_25_n_41 & {in1[13]}));
 assign mul_22_25_n_316 = ~((mul_22_25_n_60 & {in2[1]}) | (mul_22_25_n_44 & {in1[18]}));
 assign mul_22_25_n_315 = ~((mul_22_25_n_50 & {in2[11]}) | (mul_22_25_n_18 & {in1[17]}));
 assign mul_22_25_n_314 = ~((mul_22_25_n_31 & {in2[7]}) | (mul_22_25_n_20 & {in1[7]}));
 assign mul_22_25_n_313 = ~((mul_22_25_n_52 & {in2[9]}) | (mul_22_25_n_17 & {in1[6]}));
 assign mul_22_25_n_312 = ~((mul_22_25_n_50 & {in2[5]}) | (mul_22_25_n_43 & {in1[17]}));
 assign mul_22_25_n_311 = ~((mul_22_25_n_30 & {in2[9]}) | (mul_22_25_n_17 & {in1[4]}));
 assign mul_22_25_n_310 = ~((mul_22_25_n_27 & {in2[19]}) | (mul_22_25_n_41 & {in1[11]}));
 assign mul_22_25_n_309 = ~((mul_22_25_n_51 & {in2[19]}) | (mul_22_25_n_41 & {in1[16]}));
 assign mul_22_25_n_308 = ~((mul_22_25_n_61 & {in2[15]}) | (mul_22_25_n_19 & {in1[14]}));
 assign mul_22_25_n_307 = ~((mul_22_25_n_29 & {in2[17]}) | (mul_22_25_n_40 & {in1[9]}));
 assign mul_22_25_n_306 = ~((mul_22_25_n_29 & {in2[5]}) | (mul_22_25_n_43 & {in1[9]}));
 assign mul_22_25_n_304 = ~((mul_22_25_n_49 & {in2[1]}) | (mul_22_25_n_44 & {in1[12]}));
 assign mul_22_25_n_303 = ~((mul_22_25_n_27 & {in2[3]}) | (mul_22_25_n_42 & {in1[11]}));
 assign mul_22_25_n_302 = ~((mul_22_25_n_60 & {in2[9]}) | (mul_22_25_n_17 & {in1[18]}));
 assign mul_22_25_n_301 = ~((mul_22_25_n_49 & {in2[13]}) | (mul_22_25_n_21 & {in1[12]}));
 assign mul_22_25_n_300 = ~((mul_22_25_n_51 & {in2[7]}) | (mul_22_25_n_20 & {in1[16]}));
 assign mul_22_25_n_298 = ~(({in1[16]} | mul_22_25_n_44) & ({in2[1]} | mul_22_25_n_51));
 assign mul_22_25_n_297 = ~((mul_22_25_n_57 & {in2[15]}) | (mul_22_25_n_19 & {in1[5]}));
 assign mul_22_25_n_296 = ~((mul_22_25_n_49 & {in2[9]}) | (mul_22_25_n_17 & {in1[12]}));
 assign mul_22_25_n_295 = ~((mul_22_25_n_31 & {in2[11]}) | (mul_22_25_n_18 & {in1[7]}));
 assign mul_22_25_n_293 = ~((mul_22_25_n_57 & {in2[1]}) | (mul_22_25_n_44 & {in1[5]}));
 assign mul_22_25_n_292 = ~((mul_22_25_n_50 & {in2[1]}) | (mul_22_25_n_44 & {in1[17]}));
 assign mul_22_25_n_291 = ~((mul_22_25_n_28 & {in2[7]}) | (mul_22_25_n_20 & {in1[3]}));
 assign mul_22_25_n_290 = ~((mul_22_25_n_54 & {in2[19]}) | (mul_22_25_n_41 & {in1[1]}));
 assign mul_22_25_n_289 = ~((mul_22_25_n_50 & {in2[19]}) | (mul_22_25_n_41 & {in1[17]}));
 assign mul_22_25_n_288 = ~((mul_22_25_n_27 & {in2[5]}) | (mul_22_25_n_43 & {in1[11]}));
 assign mul_22_25_n_287 = ~((mul_22_25_n_57 & {in2[9]}) | (mul_22_25_n_17 & {in1[5]}));
 assign mul_22_25_n_286 = ~((mul_22_25_n_29 & {in2[3]}) | (mul_22_25_n_42 & {in1[9]}));
 assign mul_22_25_n_285 = ~((mul_22_25_n_31 & {in2[15]}) | (mul_22_25_n_19 & {in1[7]}));
 assign mul_22_25_n_284 = ~((mul_22_25_n_58 & {in2[3]}) | (mul_22_25_n_42 & {in1[8]}));
 assign mul_22_25_n_283 = ~((mul_22_25_n_48 & {in2[19]}) | (mul_22_25_n_41 & {in1[19]}));
 assign mul_22_25_n_282 = ~((mul_22_25_n_59 & {in2[3]}) | (mul_22_25_n_42 & {in1[2]}));
 assign mul_22_25_n_281 = ~((mul_22_25_n_54 & {in2[11]}) | (mul_22_25_n_18 & {in1[1]}));
 assign mul_22_25_n_280 = ~((mul_22_25_n_29 & {in2[11]}) | (mul_22_25_n_18 & {in1[9]}));
 assign mul_22_25_n_279 = ~((mul_22_25_n_53 & {in2[19]}) | (mul_22_25_n_41 & {in1[10]}));
 assign mul_22_25_n_278 = ~((mul_22_25_n_29 & {in2[9]}) | (mul_22_25_n_17 & {in1[9]}));
 assign mul_22_25_n_277 = ~((mul_22_25_n_29 & {in2[1]}) | (mul_22_25_n_44 & {in1[9]}));
 assign mul_22_25_n_276 = ~((mul_22_25_n_49 & {in2[7]}) | (mul_22_25_n_20 & {in1[12]}));
 assign mul_22_25_n_275 = ~((mul_22_25_n_49 & {in2[3]}) | (mul_22_25_n_42 & {in1[12]}));
 assign mul_22_25_n_274 = ~((mul_22_25_n_30 & {in2[3]}) | (mul_22_25_n_42 & {in1[4]}));
 assign mul_22_25_n_273 = ~((mul_22_25_n_48 & {in2[15]}) | (mul_22_25_n_19 & {in1[19]}));
 assign mul_22_25_n_272 = ~((mul_22_25_n_50 & {in2[15]}) | (mul_22_25_n_19 & {in1[17]}));
 assign mul_22_25_n_271 = ~((mul_22_25_n_59 & {in2[13]}) | (mul_22_25_n_21 & {in1[2]}));
 assign mul_22_25_n_270 = ~((mul_22_25_n_49 & {in2[19]}) | (mul_22_25_n_41 & {in1[12]}));
 assign mul_22_25_n_269 = ~((mul_22_25_n_28 & {in2[13]}) | (mul_22_25_n_21 & {in1[3]}));
 assign mul_22_25_n_268 = ~((mul_22_25_n_48 & {in2[5]}) | (mul_22_25_n_43 & {in1[19]}));
 assign mul_22_25_n_267 = ~((mul_22_25_n_30 & {in2[13]}) | (mul_22_25_n_21 & {in1[4]}));
 assign mul_22_25_n_266 = ~((mul_22_25_n_54 & {in2[15]}) | (mul_22_25_n_19 & {in1[1]}));
 assign mul_22_25_n_265 = ~((mul_22_25_n_56 & {in2[17]}) | (mul_22_25_n_40 & {in1[13]}));
 assign mul_22_25_n_264 = ~((mul_22_25_n_31 & {in2[9]}) | (mul_22_25_n_17 & {in1[7]}));
 assign mul_22_25_n_263 = ~((mul_22_25_n_48 & {in2[13]}) | (mul_22_25_n_21 & {in1[19]}));
 assign mul_22_25_n_262 = ~((mul_22_25_n_51 & {in2[11]}) | (mul_22_25_n_18 & {in1[16]}));
 assign mul_22_25_n_260 = ~((mul_22_25_n_56 & {in2[1]}) | (mul_22_25_n_44 & {in1[13]}));
 assign mul_22_25_n_259 = ~((mul_22_25_n_48 & {in2[7]}) | (mul_22_25_n_20 & {in1[19]}));
 assign mul_22_25_n_258 = ~((mul_22_25_n_52 & {in2[13]}) | (mul_22_25_n_21 & {in1[6]}));
 assign mul_22_25_n_257 = ~((mul_22_25_n_55 & {in2[9]}) | (mul_22_25_n_17 & {in1[15]}));
 assign mul_22_25_n_255 = ~(({in1[15]} | mul_22_25_n_44) & ({in2[1]} | mul_22_25_n_55));
 assign mul_22_25_n_254 = ~((mul_22_25_n_51 & {in2[5]}) | (mul_22_25_n_43 & {in1[16]}));
 assign mul_22_25_n_253 = ~((mul_22_25_n_52 & {in2[19]}) | (mul_22_25_n_41 & {in1[6]}));
 assign mul_22_25_n_252 = ~((mul_22_25_n_50 & {in2[9]}) | (mul_22_25_n_17 & {in1[17]}));
 assign mul_22_25_n_251 = ~((mul_22_25_n_58 & {in2[1]}) | (mul_22_25_n_44 & {in1[8]}));
 assign mul_22_25_n_249 = ~((mul_22_25_n_52 & {in2[1]}) | (mul_22_25_n_44 & {in1[6]}));
 assign mul_22_25_n_248 = ~((mul_22_25_n_60 & {in2[17]}) | (mul_22_25_n_40 & {in1[18]}));
 assign mul_22_25_n_247 = ~((mul_22_25_n_53 & {in2[5]}) | (mul_22_25_n_43 & {in1[10]}));
 assign mul_22_25_n_246 = ~((mul_22_25_n_53 & {in2[7]}) | (mul_22_25_n_20 & {in1[10]}));
 assign mul_22_25_n_245 = ~((mul_22_25_n_55 & {in2[15]}) | (mul_22_25_n_19 & {in1[15]}));
 assign mul_22_25_n_243 = ~(({in1[3]} | mul_22_25_n_44) & ({in2[1]} | mul_22_25_n_28));
 assign mul_22_25_n_242 = ~((mul_22_25_n_56 & {in2[9]}) | (mul_22_25_n_17 & {in1[13]}));
 assign mul_22_25_n_241 = ~((mul_22_25_n_30 & {in2[5]}) | (mul_22_25_n_43 & {in1[4]}));
 assign mul_22_25_n_239 = ~((mul_22_25_n_57 & {in2[3]}) | (mul_22_25_n_42 & {in1[5]}));
 assign mul_22_25_n_238 = ~((mul_22_25_n_30 & {in2[11]}) | (mul_22_25_n_18 & {in1[4]}));
 assign mul_22_25_n_237 = ~((mul_22_25_n_57 & {in2[5]}) | (mul_22_25_n_43 & {in1[5]}));
 assign mul_22_25_n_236 = ~((mul_22_25_n_27 & {in2[1]}) | (mul_22_25_n_44 & {in1[11]}));
 assign mul_22_25_n_234 = ~((mul_22_25_n_31 & {in2[1]}) | (mul_22_25_n_44 & {in1[7]}));
 assign mul_22_25_n_233 = ~((mul_22_25_n_31 & {in2[19]}) | (mul_22_25_n_41 & {in1[7]}));
 assign mul_22_25_n_232 = ~(({in1[2]} | mul_22_25_n_44) & ({in2[1]} | mul_22_25_n_59));
 assign mul_22_25_n_231 = ~((mul_22_25_n_59 & {in2[19]}) | (mul_22_25_n_41 & {in1[2]}));
 assign mul_22_25_n_230 = ~((mul_22_25_n_54 & {in2[13]}) | (mul_22_25_n_21 & {in1[1]}));
 assign mul_22_25_n_229 = ~((mul_22_25_n_55 & {in2[11]}) | (mul_22_25_n_18 & {in1[15]}));
 assign mul_22_25_n_228 = ~((mul_22_25_n_49 & {in2[5]}) | (mul_22_25_n_43 & {in1[12]}));
 assign mul_22_25_n_227 = ~((mul_22_25_n_56 & {in2[5]}) | (mul_22_25_n_43 & {in1[13]}));
 assign mul_22_25_n_226 = ~((mul_22_25_n_29 & {in2[7]}) | (mul_22_25_n_20 & {in1[9]}));
 assign mul_22_25_n_225 = ~((mul_22_25_n_54 & {in2[7]}) | (mul_22_25_n_20 & {in1[1]}));
 assign mul_22_25_n_224 = ~((mul_22_25_n_29 & {in2[15]}) | (mul_22_25_n_19 & {in1[9]}));
 assign mul_22_25_n_223 = ~((mul_22_25_n_33 & {in2[25]}) | (mul_22_25_n_24 & {in1[20]}));
 assign mul_22_25_n_222 = ~((mul_22_25_n_32 & {in2[25]}) | (mul_22_25_n_24 & {in1[21]}));
 assign mul_22_25_n_221 = ~((mul_22_25_n_52 & {in2[21]}) | (mul_22_25_n_22 & {in1[6]}));
 assign mul_22_25_n_220 = ~((mul_22_25_n_29 & {in2[21]}) | (mul_22_25_n_22 & {in1[9]}));
 assign mul_22_25_n_219 = ~((mul_22_25_n_58 & {in2[21]}) | (mul_22_25_n_22 & {in1[8]}));
 assign mul_22_25_n_218 = ~((mul_22_25_n_50 & {in2[21]}) | (mul_22_25_n_22 & {in1[17]}));
 assign mul_22_25_n_217 = ~((mul_22_25_n_49 & {in2[21]}) | (mul_22_25_n_22 & {in1[12]}));
 assign mul_22_25_n_216 = ~((mul_22_25_n_53 & {in2[21]}) | (mul_22_25_n_22 & {in1[10]}));
 assign mul_22_25_n_215 = ~((mul_22_25_n_27 & {in2[21]}) | (mul_22_25_n_22 & {in1[11]}));
 assign mul_22_25_n_214 = ~((mul_22_25_n_56 & {in2[21]}) | (mul_22_25_n_22 & {in1[13]}));
 assign mul_22_25_n_213 = ~((mul_22_25_n_31 & {in2[21]}) | (mul_22_25_n_22 & {in1[7]}));
 assign mul_22_25_n_212 = ~((mul_22_25_n_57 & {in2[21]}) | (mul_22_25_n_22 & {in1[5]}));
 assign mul_22_25_n_211 = ~((mul_22_25_n_59 & {in2[21]}) | (mul_22_25_n_22 & {in1[2]}));
 assign mul_22_25_n_210 = ~((mul_22_25_n_51 & {in2[21]}) | (mul_22_25_n_22 & {in1[16]}));
 assign mul_22_25_n_209 = ~((mul_22_25_n_60 & {in2[21]}) | (mul_22_25_n_22 & {in1[18]}));
 assign mul_22_25_n_208 = ~((mul_22_25_n_48 & {in2[21]}) | (mul_22_25_n_22 & {in1[19]}));
 assign mul_22_25_n_207 = ~((mul_22_25_n_54 & {in2[21]}) | (mul_22_25_n_22 & {in1[1]}));
 assign mul_22_25_n_206 = ~((mul_22_25_n_28 & {in2[21]}) | (mul_22_25_n_22 & {in1[3]}));
 assign mul_22_25_n_205 = ~((mul_22_25_n_55 & {in2[21]}) | (mul_22_25_n_22 & {in1[15]}));
 assign mul_22_25_n_204 = ~((mul_22_25_n_61 & {in2[21]}) | (mul_22_25_n_22 & {in1[14]}));
 assign mul_22_25_n_203 = ~((mul_22_25_n_30 & {in2[21]}) | (mul_22_25_n_22 & {in1[4]}));
 assign mul_22_25_n_202 = ~((mul_22_25_n_29 & {in2[23]}) | (mul_22_25_n_45 & {in1[9]}));
 assign mul_22_25_n_201 = ~((mul_22_25_n_56 & {in2[23]}) | (mul_22_25_n_45 & {in1[13]}));
 assign mul_22_25_n_200 = ~((mul_22_25_n_54 & {in2[23]}) | (mul_22_25_n_45 & {in1[1]}));
 assign mul_22_25_n_199 = ~((mul_22_25_n_30 & {in2[23]}) | (mul_22_25_n_45 & {in1[4]}));
 assign mul_22_25_n_198 = ~((mul_22_25_n_53 & {in2[23]}) | (mul_22_25_n_45 & {in1[10]}));
 assign mul_22_25_n_197 = ~((mul_22_25_n_61 & {in2[23]}) | (mul_22_25_n_45 & {in1[14]}));
 assign mul_22_25_n_196 = ~((mul_22_25_n_49 & {in2[23]}) | (mul_22_25_n_45 & {in1[12]}));
 assign mul_22_25_n_195 = ~((mul_22_25_n_31 & {in2[23]}) | (mul_22_25_n_45 & {in1[7]}));
 assign mul_22_25_n_194 = ~((mul_22_25_n_55 & {in2[23]}) | (mul_22_25_n_45 & {in1[15]}));
 assign mul_22_25_n_193 = ~((mul_22_25_n_27 & {in2[23]}) | (mul_22_25_n_45 & {in1[11]}));
 assign mul_22_25_n_192 = ~((mul_22_25_n_58 & {in2[23]}) | (mul_22_25_n_45 & {in1[8]}));
 assign mul_22_25_n_191 = ~((mul_22_25_n_50 & {in2[23]}) | (mul_22_25_n_45 & {in1[17]}));
 assign mul_22_25_n_190 = ~((mul_22_25_n_57 & {in2[23]}) | (mul_22_25_n_45 & {in1[5]}));
 assign mul_22_25_n_189 = ~((mul_22_25_n_51 & {in2[23]}) | (mul_22_25_n_45 & {in1[16]}));
 assign mul_22_25_n_188 = ~((mul_22_25_n_60 & {in2[23]}) | (mul_22_25_n_45 & {in1[18]}));
 assign mul_22_25_n_187 = ~((mul_22_25_n_52 & {in2[23]}) | (mul_22_25_n_45 & {in1[6]}));
 assign mul_22_25_n_186 = ~((mul_22_25_n_28 & {in2[23]}) | (mul_22_25_n_45 & {in1[3]}));
 assign mul_22_25_n_185 = ~((mul_22_25_n_59 & {in2[23]}) | (mul_22_25_n_45 & {in1[2]}));
 assign mul_22_25_n_184 = ~((mul_22_25_n_48 & {in2[23]}) | (mul_22_25_n_45 & {in1[19]}));
 assign mul_22_25_n_183 = ~((mul_22_25_n_32 & {in2[27]}) | (mul_22_25_n_25 & {in1[21]}));
 assign mul_22_25_n_182 = ~((mul_22_25_n_33 & {in2[27]}) | (mul_22_25_n_25 & {in1[20]}));
 assign mul_22_25_n_181 = ~((mul_22_25_n_51 & {in2[3]}) | (mul_22_25_n_42 & {in1[16]}));
 assign mul_22_25_n_180 = ~((mul_22_25_n_30 & {in2[25]}) | (mul_22_25_n_24 & {in1[4]}));
 assign mul_22_25_n_179 = ~((mul_22_25_n_31 & {in2[25]}) | (mul_22_25_n_24 & {in1[7]}));
 assign mul_22_25_n_178 = ~((mul_22_25_n_27 & {in2[25]}) | (mul_22_25_n_24 & {in1[11]}));
 assign mul_22_25_n_177 = ~((mul_22_25_n_56 & {in2[25]}) | (mul_22_25_n_24 & {in1[13]}));
 assign mul_22_25_n_176 = ~((mul_22_25_n_29 & {in2[25]}) | (mul_22_25_n_24 & {in1[9]}));
 assign mul_22_25_n_175 = ~((mul_22_25_n_52 & {in2[25]}) | (mul_22_25_n_24 & {in1[6]}));
 assign mul_22_25_n_174 = ~((mul_22_25_n_57 & {in2[25]}) | (mul_22_25_n_24 & {in1[5]}));
 assign mul_22_25_n_173 = ~((mul_22_25_n_54 & {in2[25]}) | (mul_22_25_n_24 & {in1[1]}));
 assign mul_22_25_n_172 = ~((mul_22_25_n_58 & {in2[25]}) | (mul_22_25_n_24 & {in1[8]}));
 assign mul_22_25_n_171 = ~((mul_22_25_n_61 & {in2[25]}) | (mul_22_25_n_24 & {in1[14]}));
 assign mul_22_25_n_170 = ~((mul_22_25_n_28 & {in2[25]}) | (mul_22_25_n_24 & {in1[3]}));
 assign mul_22_25_n_169 = ~((mul_22_25_n_51 & {in2[25]}) | (mul_22_25_n_24 & {in1[16]}));
 assign mul_22_25_n_168 = ~((mul_22_25_n_48 & {in2[25]}) | (mul_22_25_n_24 & {in1[19]}));
 assign mul_22_25_n_167 = ~((mul_22_25_n_53 & {in2[25]}) | (mul_22_25_n_24 & {in1[10]}));
 assign mul_22_25_n_166 = ~((mul_22_25_n_59 & {in2[25]}) | (mul_22_25_n_24 & {in1[2]}));
 assign mul_22_25_n_165 = ~((mul_22_25_n_60 & {in2[25]}) | (mul_22_25_n_24 & {in1[18]}));
 assign mul_22_25_n_164 = ~((mul_22_25_n_55 & {in2[25]}) | (mul_22_25_n_24 & {in1[15]}));
 assign mul_22_25_n_163 = ~((mul_22_25_n_49 & {in2[25]}) | (mul_22_25_n_24 & {in1[12]}));
 assign mul_22_25_n_162 = ~((mul_22_25_n_50 & {in2[25]}) | (mul_22_25_n_24 & {in1[17]}));
 assign mul_22_25_n_161 = ~((mul_22_25_n_33 & {in2[29]}) | (mul_22_25_n_46 & {in1[20]}));
 assign mul_22_25_n_160 = ~((mul_22_25_n_53 & {in2[9]}) | (mul_22_25_n_17 & {in1[10]}));
 assign mul_22_25_n_159 = ~((mul_22_25_n_48 & {in2[27]}) | (mul_22_25_n_25 & {in1[19]}));
 assign mul_22_25_n_158 = ~((mul_22_25_n_56 & {in2[27]}) | (mul_22_25_n_25 & {in1[13]}));
 assign mul_22_25_n_157 = ~((mul_22_25_n_61 & {in2[27]}) | (mul_22_25_n_25 & {in1[14]}));
 assign mul_22_25_n_156 = ~((mul_22_25_n_54 & {in2[27]}) | (mul_22_25_n_25 & {in1[1]}));
 assign mul_22_25_n_155 = ~((mul_22_25_n_30 & {in2[27]}) | (mul_22_25_n_25 & {in1[4]}));
 assign mul_22_25_n_154 = ~((mul_22_25_n_27 & {in2[27]}) | (mul_22_25_n_25 & {in1[11]}));
 assign mul_22_25_n_153 = ~((mul_22_25_n_29 & {in2[27]}) | (mul_22_25_n_25 & {in1[9]}));
 assign mul_22_25_n_152 = ~((mul_22_25_n_53 & {in2[27]}) | (mul_22_25_n_25 & {in1[10]}));
 assign mul_22_25_n_151 = ~((mul_22_25_n_59 & {in2[27]}) | (mul_22_25_n_25 & {in1[2]}));
 assign mul_22_25_n_150 = ~((mul_22_25_n_28 & {in2[27]}) | (mul_22_25_n_25 & {in1[3]}));
 assign mul_22_25_n_149 = ~((mul_22_25_n_51 & {in2[27]}) | (mul_22_25_n_25 & {in1[16]}));
 assign mul_22_25_n_148 = ~((mul_22_25_n_58 & {in2[27]}) | (mul_22_25_n_25 & {in1[8]}));
 assign mul_22_25_n_147 = ~((mul_22_25_n_31 & {in2[27]}) | (mul_22_25_n_25 & {in1[7]}));
 assign mul_22_25_n_146 = ~((mul_22_25_n_55 & {in2[27]}) | (mul_22_25_n_25 & {in1[15]}));
 assign mul_22_25_n_145 = ~((mul_22_25_n_60 & {in2[27]}) | (mul_22_25_n_25 & {in1[18]}));
 assign mul_22_25_n_144 = ~((mul_22_25_n_52 & {in2[27]}) | (mul_22_25_n_25 & {in1[6]}));
 assign mul_22_25_n_143 = ~((mul_22_25_n_57 & {in2[27]}) | (mul_22_25_n_25 & {in1[5]}));
 assign mul_22_25_n_142 = ~((mul_22_25_n_49 & {in2[27]}) | (mul_22_25_n_25 & {in1[12]}));
 assign mul_22_25_n_141 = ~((mul_22_25_n_50 & {in2[27]}) | (mul_22_25_n_25 & {in1[17]}));
 assign mul_22_25_n_140 = ~((mul_22_25_n_29 & {in2[29]}) | (mul_22_25_n_46 & {in1[9]}));
 assign mul_22_25_n_139 = ~((mul_22_25_n_55 & {in2[29]}) | (mul_22_25_n_46 & {in1[15]}));
 assign mul_22_25_n_138 = ~((mul_22_25_n_57 & {in2[29]}) | (mul_22_25_n_46 & {in1[5]}));
 assign mul_22_25_n_137 = ~((mul_22_25_n_48 & {in2[29]}) | (mul_22_25_n_46 & {in1[19]}));
 assign mul_22_25_n_136 = ~((mul_22_25_n_58 & {in2[29]}) | (mul_22_25_n_46 & {in1[8]}));
 assign mul_22_25_n_135 = ~((mul_22_25_n_51 & {in2[29]}) | (mul_22_25_n_46 & {in1[16]}));
 assign mul_22_25_n_134 = ~((mul_22_25_n_28 & {in2[29]}) | (mul_22_25_n_46 & {in1[3]}));
 assign mul_22_25_n_133 = ~((mul_22_25_n_50 & {in2[29]}) | (mul_22_25_n_46 & {in1[17]}));
 assign mul_22_25_n_132 = ~((mul_22_25_n_54 & {in2[29]}) | (mul_22_25_n_46 & {in1[1]}));
 assign mul_22_25_n_131 = ~((mul_22_25_n_30 & {in2[29]}) | (mul_22_25_n_46 & {in1[4]}));
 assign mul_22_25_n_130 = ~((mul_22_25_n_60 & {in2[29]}) | (mul_22_25_n_46 & {in1[18]}));
 assign mul_22_25_n_129 = ~((mul_22_25_n_56 & {in2[29]}) | (mul_22_25_n_46 & {in1[13]}));
 assign mul_22_25_n_128 = ~((mul_22_25_n_31 & {in2[29]}) | (mul_22_25_n_46 & {in1[7]}));
 assign mul_22_25_n_127 = ~((mul_22_25_n_27 & {in2[29]}) | (mul_22_25_n_46 & {in1[11]}));
 assign mul_22_25_n_126 = ~((mul_22_25_n_53 & {in2[29]}) | (mul_22_25_n_46 & {in1[10]}));
 assign mul_22_25_n_125 = ~((mul_22_25_n_49 & {in2[29]}) | (mul_22_25_n_46 & {in1[12]}));
 assign mul_22_25_n_124 = ~((mul_22_25_n_59 & {in2[29]}) | (mul_22_25_n_46 & {in1[2]}));
 assign mul_22_25_n_123 = ~((mul_22_25_n_52 & {in2[29]}) | (mul_22_25_n_46 & {in1[6]}));
 assign mul_22_25_n_122 = ~((mul_22_25_n_61 & {in2[29]}) | (mul_22_25_n_46 & {in1[14]}));
 assign mul_22_25_n_121 = ~((mul_22_25_n_27 & {in2[31]}) | (mul_22_25_n_47 & {in1[11]}));
 assign mul_22_25_n_120 = ~((mul_22_25_n_60 & {in2[31]}) | (mul_22_25_n_47 & {in1[18]}));
 assign mul_22_25_n_119 = ~((mul_22_25_n_53 & {in2[31]}) | (mul_22_25_n_47 & {in1[10]}));
 assign mul_22_25_n_118 = ~((mul_22_25_n_31 & {in2[31]}) | (mul_22_25_n_47 & {in1[7]}));
 assign mul_22_25_n_117 = ~((mul_22_25_n_61 & {in2[31]}) | (mul_22_25_n_47 & {in1[14]}));
 assign mul_22_25_n_116 = ~((mul_22_25_n_52 & {in2[31]}) | (mul_22_25_n_47 & {in1[6]}));
 assign mul_22_25_n_115 = ~((mul_22_25_n_55 & {in2[19]}) | (mul_22_25_n_41 & {in1[15]}));
 assign mul_22_25_n_114 = ~((mul_22_25_n_56 & {in2[31]}) | (mul_22_25_n_47 & {in1[13]}));
 assign mul_22_25_n_113 = ~((mul_22_25_n_55 & {in2[31]}) | (mul_22_25_n_47 & {in1[15]}));
 assign mul_22_25_n_112 = ~((mul_22_25_n_30 & {in2[31]}) | (mul_22_25_n_47 & {in1[4]}));
 assign mul_22_25_n_111 = ~((mul_22_25_n_50 & {in2[31]}) | (mul_22_25_n_47 & {in1[17]}));
 assign mul_22_25_n_110 = ~((mul_22_25_n_29 & {in2[31]}) | (mul_22_25_n_47 & {in1[9]}));
 assign mul_22_25_n_109 = ~((mul_22_25_n_51 & {in2[31]}) | (mul_22_25_n_47 & {in1[16]}));
 assign mul_22_25_n_108 = ~((mul_22_25_n_54 & {in2[31]}) | (mul_22_25_n_47 & {in1[1]}));
 assign mul_22_25_n_107 = ~((mul_22_25_n_49 & {in2[31]}) | (mul_22_25_n_47 & {in1[12]}));
 assign mul_22_25_n_106 = ~((mul_22_25_n_59 & {in2[31]}) | (mul_22_25_n_47 & {in1[2]}));
 assign mul_22_25_n_105 = ~((mul_22_25_n_28 & {in2[31]}) | (mul_22_25_n_47 & {in1[3]}));
 assign mul_22_25_n_104 = ~((mul_22_25_n_57 & {in2[31]}) | (mul_22_25_n_47 & {in1[5]}));
 assign mul_22_25_n_103 = ~((mul_22_25_n_58 & {in2[31]}) | (mul_22_25_n_47 & {in1[8]}));
 assign mul_22_25_n_102 = ~((mul_22_25_n_53 & {in2[13]}) | (mul_22_25_n_21 & {in1[10]}));
 assign mul_22_25_n_101 = ~((mul_22_25_n_27 & {in2[15]}) | (mul_22_25_n_19 & {in1[11]}));
 assign mul_22_25_n_100 = ~((mul_22_25_n_61 & {in2[3]}) | (mul_22_25_n_42 & {in1[14]}));
 assign mul_22_25_n_99 = ~((mul_22_25_n_56 & {in2[7]}) | (mul_22_25_n_20 & {in1[13]}));
 assign mul_22_25_n_98 = ~((mul_22_25_n_52 & {in2[11]}) | (mul_22_25_n_18 & {in1[6]}));
 assign mul_22_25_n_97 = ~((mul_22_25_n_60 & {in2[5]}) | (mul_22_25_n_43 & {in1[18]}));
 assign mul_22_25_n_96 = ~((mul_22_25_n_50 & {in2[3]}) | (mul_22_25_n_42 & {in1[17]}));
 assign mul_22_25_n_95 = ~((mul_22_25_n_28 & {in2[9]}) | (mul_22_25_n_17 & {in1[3]}));
 assign mul_22_25_n_94 = ~((mul_22_25_n_27 & {in2[11]}) | (mul_22_25_n_18 & {in1[11]}));
 assign mul_22_25_n_92 = ~(({in1[4]} | mul_22_25_n_44) & ({in2[1]} | mul_22_25_n_30));
 assign mul_22_25_n_91 = ~((mul_22_25_n_52 & {in2[17]}) | (mul_22_25_n_40 & {in1[6]}));
 assign mul_22_25_n_90 = ~((mul_22_25_n_59 & {in2[15]}) | (mul_22_25_n_19 & {in1[2]}));
 assign mul_22_25_n_89 = ~((mul_22_25_n_59 & {in2[7]}) | (mul_22_25_n_20 & {in1[2]}));
 assign mul_22_25_n_88 = ~((mul_22_25_n_58 & {in2[15]}) | (mul_22_25_n_19 & {in1[8]}));
 assign mul_22_25_n_87 = ~((mul_22_25_n_50 & {in2[7]}) | (mul_22_25_n_20 & {in1[17]}));
 assign mul_22_25_n_86 = ~((mul_22_25_n_50 & {in2[17]}) | (mul_22_25_n_40 & {in1[17]}));
 assign asc001_0_ = ~(mul_22_25_n_26 | mul_22_25_n_23);
 assign mul_22_25_n_65 = ~{in1[29]};
 assign mul_22_25_n_64 = ~{in1[28]};
 assign mul_22_25_n_63 = ~{in1[27]};
 assign mul_22_25_n_62 = ~{in1[25]};
 assign mul_22_25_n_61 = ~{in1[14]};
 assign mul_22_25_n_60 = ~{in1[18]};
 assign mul_22_25_n_59 = ~{in1[2]};
 assign mul_22_25_n_58 = ~{in1[8]};
 assign mul_22_25_n_57 = ~{in1[5]};
 assign mul_22_25_n_56 = ~{in1[13]};
 assign mul_22_25_n_55 = ~{in1[15]};
 assign mul_22_25_n_54 = ~{in1[1]};
 assign mul_22_25_n_53 = ~{in1[10]};
 assign mul_22_25_n_52 = ~{in1[6]};
 assign mul_22_25_n_51 = ~{in1[16]};
 assign mul_22_25_n_50 = ~{in1[17]};
 assign mul_22_25_n_49 = ~{in1[12]};
 assign mul_22_25_n_48 = ~{in1[19]};
 assign mul_22_25_n_47 = ~{in2[31]};
 assign mul_22_25_n_46 = ~{in2[29]};
 assign mul_22_25_n_45 = ~{in2[23]};
 assign mul_22_25_n_44 = ~{in2[1]};
 assign mul_22_25_n_43 = ~{in2[5]};
 assign mul_22_25_n_42 = ~{in2[3]};
 assign mul_22_25_n_41 = ~{in2[19]};
 assign mul_22_25_n_40 = ~{in2[17]};
 assign mul_22_25_n_39 = ~{in1[30]};
 assign mul_22_25_n_38 = ~{in1[31]};
 assign mul_22_25_n_37 = ~{in1[26]};
 assign mul_22_25_n_36 = ~{in1[24]};
 assign mul_22_25_n_35 = ~{in1[22]};
 assign mul_22_25_n_34 = ~{in1[23]};
 assign mul_22_25_n_33 = ~{in1[20]};
 assign mul_22_25_n_32 = ~{in1[21]};
 assign mul_22_25_n_31 = ~{in1[7]};
 assign mul_22_25_n_30 = ~{in1[4]};
 assign mul_22_25_n_29 = ~{in1[9]};
 assign mul_22_25_n_28 = ~{in1[3]};
 assign mul_22_25_n_27 = ~{in1[11]};
 assign mul_22_25_n_26 = ~{in2[0]};
 assign mul_22_25_n_25 = ~{in2[27]};
 assign mul_22_25_n_24 = ~{in2[25]};
 assign mul_22_25_n_23 = ~{in1[0]};
 assign mul_22_25_n_22 = ~{in2[21]};
 assign mul_22_25_n_21 = ~{in2[13]};
 assign mul_22_25_n_20 = ~{in2[7]};
 assign mul_22_25_n_19 = ~{in2[15]};
 assign mul_22_25_n_18 = ~{in2[11]};
 assign mul_22_25_n_17 = ~{in2[9]};
 assign mul_22_25_n_15 = (mul_22_25_n_2244 | mul_22_25_n_2283);
 assign asc001_22_ = (mul_22_25_n_1338 ^ mul_22_25_n_1376);
 assign mul_22_25_n_13 = ~(mul_22_25_n_1314 | (~mul_22_25_n_1375 & mul_22_25_n_1312));
 assign mul_22_25_n_12 = (mul_22_25_n_2251 | mul_22_25_n_2290);
 assign mul_22_25_n_11 = ~(mul_22_25_n_1302 & (~mul_22_25_n_1366 | mul_22_25_n_1305));
 assign mul_22_25_n_10 = (mul_22_25_n_2264 ^ n_137);
 assign mul_22_25_n_9 = (n_96 | n_135);
 assign asc001_10_ = ~(mul_22_25_n_1228 ^ mul_22_25_n_1236);
 assign mul_22_25_n_7 = ~(~mul_22_25_n_355 & mul_22_25_n_566);
 assign mul_22_25_n_6 = ~(~mul_22_25_n_357 & mul_22_25_n_565);
 assign mul_22_25_n_5 = ~(~mul_22_25_n_356 & mul_22_25_n_570);
 assign mul_22_25_n_4 = ~(~mul_22_25_n_352 & mul_22_25_n_572);
 assign mul_22_25_n_3 = ~(~mul_22_25_n_350 & mul_22_25_n_567);
 assign mul_22_25_n_2 = ~(mul_22_25_n_353 | ~mul_22_25_n_575);
 assign mul_22_25_n_1 = ~(mul_22_25_n_640 | (~mul_22_25_n_573 & mul_22_25_n_601));
 assign mul_22_25_n_0 = ~(mul_22_25_n_2 | (~mul_22_25_n_563 & mul_22_25_n_609));
 assign n_0 = ~clr;
 assign mul_22_25_n_1535 = (mul_22_25_n_1072 ^ (mul_22_25_n_1073 ^ mul_22_25_n_1076));
 assign mul_22_25_n_1534 = (mul_22_25_n_1074 ^ (mul_22_25_n_1075 ^ mul_22_25_n_1077));
 assign mul_22_25_n_1532 = (mul_22_25_n_1536 ^ (mul_22_25_n_1537 ^ mul_22_25_n_1078));
 assign mul_22_25_n_1530 = (mul_22_25_n_1533 ^ (mul_22_25_n_1534 ^ mul_22_25_n_1535));
 assign mul_22_25_n_1528 = (mul_22_25_n_1530 ^ (mul_22_25_n_1531 ^ mul_22_25_n_1532));
 assign mul_22_25_n_2303 = (mul_22_25_n_1527 ^ (mul_22_25_n_1528 ^ mul_22_25_n_1529));
endmodule


