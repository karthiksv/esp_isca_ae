`timescale 1ps / 1ps
module divider_hls_Div_13Ux7U_6U_4(
          in2,
          in1,
          out1,
          clk,
          rst
);
   input [12:0] in2;
   input [6:0] in1;
   output [5:0] out1;
   input clk;
   input rst;
wire rst, clk, n_51, n_52, n_53, n_54, n_55, n_56, n_148, n_149, n_150, n_151,
     n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_162, n_163,
     n_164, n_165, n_167, n_168, n_169, n_171, n_172, n_173, n_180, n_181, n_182,
     n_183, n_184, n_185, n_186, n_25, n_26, n_27, sub_149_2_n_1, sub_149_2_n_2,
     sub_149_2_n_3, sub_149_2_n_4, sub_149_2_n_5, sub_149_2_n_6, sub_149_2_n_7,
     sub_149_2_n_8, sub_149_2_n_9, sub_149_2_n_10, sub_149_2_n_11,
     sub_149_2_n_12, sub_149_2_n_13, sub_149_2_n_14, sub_149_2_n_15,
     sub_149_2_n_16, sub_149_2_n_17, sub_149_2_n_19, sub_149_2_n_20,
     sub_149_2_n_21, sub_149_2_n_22, sub_149_2_n_23, sub_149_2_n_24,
     sub_149_2_n_25, sub_149_2_n_26, sub_149_2_n_27, sub_149_2_n_29,
     sub_149_2_n_30, sub_149_2_n_32, sub_149_2_n_33, sub_248_2_n_0,
     sub_248_2_n_1, sub_248_2_n_2, sub_248_2_n_3, sub_248_2_n_4, sub_248_2_n_5,
     sub_248_2_n_6, sub_248_2_n_7, sub_248_2_n_8, sub_248_2_n_9, sub_248_2_n_10,
     sub_248_2_n_11, sub_248_2_n_12, sub_248_2_n_13, sub_248_2_n_14,
     sub_248_2_n_15, sub_248_2_n_16, sub_248_2_n_18, sub_248_2_n_19,
     sub_248_2_n_20, sub_248_2_n_21, sub_248_2_n_22, sub_248_2_n_23,
     sub_248_2_n_24, sub_248_2_n_25, sub_248_2_n_26, sub_248_2_n_27,
     sub_248_2_n_28, sub_248_2_n_30, sub_248_2_n_32, sub_248_2_n_33,
     sub_248_2_n_34, sub_248_2_n_35, sub_248_2_n_36, sub_248_2_n_39,
     sub_248_2_n_40, sub_248_2_n_41, sub_168_2_n_0, sub_168_2_n_1, sub_168_2_n_2,
     sub_168_2_n_3, sub_168_2_n_4, sub_168_2_n_5, sub_168_2_n_6, sub_168_2_n_7,
     sub_168_2_n_8, sub_168_2_n_9, sub_168_2_n_10, sub_168_2_n_11,
     sub_168_2_n_12, sub_168_2_n_13, sub_168_2_n_14, sub_168_2_n_15,
     sub_168_2_n_16, sub_168_2_n_17, sub_168_2_n_18, sub_168_2_n_20,
     sub_168_2_n_21, sub_168_2_n_22, sub_168_2_n_23, sub_168_2_n_24,
     sub_168_2_n_25, sub_168_2_n_26, sub_168_2_n_27, sub_168_2_n_28,
     sub_168_2_n_29, sub_168_2_n_30, sub_168_2_n_32, sub_168_2_n_33,
     sub_168_2_n_34, sub_168_2_n_36, sub_168_2_n_37, sub_168_2_n_38,
     sub_168_2_n_39, sub_168_2_n_40, sub_168_2_n_43, sub_187_2_n_0,
     sub_187_2_n_1, sub_187_2_n_2, sub_187_2_n_3, sub_187_2_n_4, sub_187_2_n_5,
     sub_187_2_n_6, sub_187_2_n_7, sub_187_2_n_8, sub_187_2_n_9, sub_187_2_n_10,
     sub_187_2_n_11, sub_187_2_n_12, sub_187_2_n_13, sub_187_2_n_14,
     sub_187_2_n_15, sub_187_2_n_16, sub_187_2_n_17, sub_187_2_n_18,
     sub_187_2_n_19, sub_187_2_n_20, sub_187_2_n_21, sub_187_2_n_22,
     sub_187_2_n_23, sub_187_2_n_24, sub_187_2_n_25, sub_187_2_n_26,
     sub_187_2_n_27, sub_187_2_n_29, sub_187_2_n_30, sub_187_2_n_31,
     sub_187_2_n_32, sub_187_2_n_33, sub_187_2_n_34, sub_187_2_n_35,
     sub_187_2_n_36, sub_187_2_n_37, sub_187_2_n_38, sub_187_2_n_39,
     sub_187_2_n_41, sub_187_2_n_42, sub_187_2_n_43, sub_187_2_n_45,
     sub_187_2_n_46, sub_187_2_n_47, sub_187_2_n_48, sub_187_2_n_49,
     sub_187_2_n_50, sub_187_2_n_51, sub_187_2_n_54, sub_187_2_n_55,
     sub_269_2_n_0, sub_269_2_n_1, sub_269_2_n_2, sub_269_2_n_3, sub_269_2_n_4,
     sub_269_2_n_5, sub_269_2_n_6, sub_269_2_n_7, sub_269_2_n_8, sub_269_2_n_9,
     sub_269_2_n_10, sub_269_2_n_11, sub_269_2_n_12, sub_269_2_n_13,
     sub_269_2_n_14, sub_269_2_n_15, sub_269_2_n_16, sub_269_2_n_18,
     sub_269_2_n_19, sub_269_2_n_20, sub_269_2_n_21, sub_269_2_n_22,
     sub_269_2_n_23, sub_269_2_n_24, sub_269_2_n_25, sub_269_2_n_26,
     sub_269_2_n_27, sub_269_2_n_28, sub_269_2_n_30, sub_269_2_n_32,
     sub_269_2_n_33, sub_269_2_n_34, sub_269_2_n_35, sub_269_2_n_36,
     sub_269_2_n_39, sub_269_2_n_40, sub_269_2_n_41, sub_290_2_n_0,
     sub_290_2_n_1, sub_290_2_n_2, sub_290_2_n_3, sub_290_2_n_4, sub_290_2_n_5,
     sub_290_2_n_6, sub_290_2_n_7, sub_290_2_n_8, sub_290_2_n_9, sub_290_2_n_10,
     sub_290_2_n_11, sub_290_2_n_12, sub_290_2_n_13, sub_290_2_n_14,
     sub_290_2_n_15, sub_290_2_n_16, sub_290_2_n_18, sub_290_2_n_19,
     sub_290_2_n_20, sub_290_2_n_21, sub_290_2_n_22, sub_290_2_n_23,
     sub_290_2_n_24, sub_290_2_n_25, sub_290_2_n_26, sub_290_2_n_27,
     sub_290_2_n_28, sub_290_2_n_30, sub_290_2_n_32, sub_290_2_n_33,
     sub_290_2_n_34, sub_290_2_n_35, sub_290_2_n_36, sub_290_2_n_39,
     sub_290_2_n_40, sub_290_2_n_41, sub_206_2_n_0, sub_206_2_n_1, sub_206_2_n_2,
     sub_206_2_n_3, sub_206_2_n_6, sub_206_2_n_7, sub_206_2_n_8, sub_206_2_n_9,
     sub_206_2_n_10, sub_206_2_n_11, sub_206_2_n_12, sub_206_2_n_13,
     sub_206_2_n_14, sub_206_2_n_15, sub_206_2_n_16, sub_206_2_n_17,
     sub_206_2_n_18, sub_206_2_n_19, sub_206_2_n_21, sub_206_2_n_22,
     sub_206_2_n_24, sub_206_2_n_25, sub_206_2_n_26, sub_206_2_n_27,
     sub_206_2_n_28, sub_206_2_n_29, sub_206_2_n_30, sub_206_2_n_31,
     sub_206_2_n_32, sub_206_2_n_33, sub_206_2_n_35, sub_206_2_n_36,
     sub_206_2_n_37, sub_206_2_n_39, sub_206_2_n_40, sub_206_2_n_41,
     sub_206_2_n_42, sub_206_2_n_43, sub_206_2_n_44, sub_206_2_n_47,
     sub_206_2_n_48, sub_206_2_n_49, sub_206_2_n_77, sub_206_2_n_78,
     sub_206_2_n_79, sub_206_2_n_81, sub_206_2_n_82, sub_206_2_n_83,
     sub_206_2_n_84, sub_206_2_n_85, sub_73_2_n_1, sub_73_2_n_2, sub_73_2_n_4,
     sub_73_2_n_5, sub_73_2_n_6, sub_92_2_n_1, sub_92_2_n_2, sub_92_2_n_3,
     sub_92_2_n_4, sub_92_2_n_5, sub_92_2_n_6, sub_92_2_n_8, sub_92_2_n_9,
     sub_111_2_n_1, sub_111_2_n_2, sub_111_2_n_3, sub_111_2_n_4, sub_111_2_n_5,
     sub_111_2_n_6, sub_111_2_n_7, sub_111_2_n_8, sub_111_2_n_10, sub_111_2_n_11,
     sub_111_2_n_12, sub_111_2_n_13, sub_111_2_n_16, sub_111_2_n_17,
     sub_227_2_n_0, sub_227_2_n_1, sub_227_2_n_2, sub_227_2_n_3, sub_227_2_n_4,
     sub_227_2_n_5, sub_227_2_n_6, sub_227_2_n_7, sub_227_2_n_8, sub_227_2_n_9,
     sub_227_2_n_10, sub_227_2_n_11, sub_227_2_n_12, sub_227_2_n_13,
     sub_227_2_n_14, sub_227_2_n_15, sub_227_2_n_16, sub_227_2_n_18,
     sub_227_2_n_19, sub_227_2_n_20, sub_227_2_n_21, sub_227_2_n_22,
     sub_227_2_n_23, sub_227_2_n_24, sub_227_2_n_25, sub_227_2_n_26,
     sub_227_2_n_27, sub_227_2_n_28, sub_227_2_n_30, sub_227_2_n_32,
     sub_227_2_n_33, sub_227_2_n_34, sub_227_2_n_35, sub_227_2_n_36,
     sub_227_2_n_39, sub_227_2_n_40, sub_227_2_n_41, sub_309_2_n_1,
     sub_309_2_n_2, sub_309_2_n_3, sub_309_2_n_4, sub_309_2_n_5, sub_309_2_n_6,
     sub_309_2_n_7, sub_309_2_n_8, sub_309_2_n_9, sub_309_2_n_10, sub_309_2_n_12,
     sub_309_2_n_13, sub_309_2_n_14, sub_309_2_n_15, sub_309_2_n_16,
     sub_309_2_n_17, sub_309_2_n_18, sub_309_2_n_19, sub_309_2_n_20,
     sub_309_2_n_21, sub_309_2_n_22, sub_309_2_n_23, sub_309_2_n_24,
     sub_309_2_n_25, sub_309_2_n_0, sub_309_2_n_47, sub_130_2_n_1, sub_130_2_n_2,
     sub_130_2_n_3, sub_130_2_n_4, sub_130_2_n_5, sub_130_2_n_6, sub_130_2_n_7,
     sub_130_2_n_8, sub_130_2_n_9, sub_130_2_n_10, sub_130_2_n_11,
     sub_130_2_n_13, sub_130_2_n_14, sub_130_2_n_15, sub_130_2_n_16,
     sub_130_2_n_17, sub_130_2_n_18, sub_130_2_n_19, sub_130_2_n_20,
     sub_130_2_n_22, sub_130_2_n_23, sub_130_2_n_25, sub_130_2_n_26,
     sub_130_2_n_27, asc001_0_0_, asc001_0_1_, asc001_0_2_, asc001_0_3_,
     asc001_0_4_, asc001_0_5_, in2_1_0_, in2_1_7_, in2_2_0_, in2_4_0_, in2_4_1_,
     in2_4_7_, in2_5_0_, in2_5_1_, in2_7_0_, in2_7_1_, in2_7_2_, in2_7_7_,
     in2_8_0_, in2_8_1_, in2_8_2_, in2_10_0_, in2_10_1_, in2_10_2_, in2_10_3_,
     in2_10_7_, in2_11_0_, in2_11_1_, in2_11_2_, in2_11_3_, in2_13_0_, in2_13_1_,
     in2_13_2_, in2_13_3_, in2_13_4_, in2_13_7_, in2_14_0_, in2_14_1_, in2_14_2_,
     in2_14_3_, in2_14_4_, in2_16_0_, in2_16_1_, in2_16_2_, in2_16_3_, in2_16_4_,
     in2_16_5_, in2_16_7_, in2_17_0_, in2_17_1_, in2_17_2_, in2_17_3_, in2_17_4_,
     in2_17_5_, in2_19_0_, in2_19_1_, in2_19_2_, in2_19_3_, in2_19_4_, in2_19_5_,
     in2_19_6_, in2_19_7_, in2_20_6_, in2_22_0_, in2_22_1_, in2_22_2_, in2_22_3_,
     in2_22_4_, in2_22_5_, in2_22_6_, in2_22_7_, in2_23_0_, in2_23_1_, in2_23_2_,
     in2_23_3_, in2_23_4_, in2_23_5_, in2_23_6_, in2_25_0_, in2_25_1_, in2_25_2_,
     in2_25_3_, in2_25_4_, in2_25_5_, in2_25_6_, in2_25_7_, in2_26_0_, in2_26_1_,
     in2_26_2_, in2_26_3_, in2_26_4_, in2_26_5_, in2_26_6_, in2_28_0_, in2_28_1_,
     in2_28_2_, in2_28_3_, in2_28_4_, in2_28_5_, in2_28_6_, in2_28_7_, in2_29_0_,
     in2_29_1_, in2_29_2_, in2_29_3_, in2_29_4_, in2_29_5_, in2_29_6_, in2_31_0_,
     in2_31_1_, in2_31_2_, in2_31_3_, in2_31_4_, in2_31_5_, in2_31_6_, in2_31_7_,
     in2_32_0_, in2_32_1_, in2_32_2_, in2_32_3_, in2_32_4_, in2_32_5_, in2_32_6_,
     in2_34_0_, in2_34_1_, in2_34_2_, in2_34_3_, in2_34_4_, in2_34_5_, in2_34_6_,
     in2_34_7_, in2_35_0_, in2_35_1_, in2_35_2_, in2_35_3_, in2_35_4_, in2_35_5_,
     in2_35_6_, in2_37_7_;
assign {out1[5]} = n_51;
assign {out1[4]} = n_52;
assign {out1[3]} = n_53;
assign {out1[2]} = n_54;
assign {out1[1]} = n_55;
assign {out1[0]} = n_56;
 reg retime_s1_2_reg_reg_IQ;
 always @(posedge clk)
         retime_s1_2_reg_reg_IQ <= n_186;
 assign n_155 = retime_s1_2_reg_reg_IQ;
 reg retime_s1_6_reg_reg_IQ;
 always @(posedge clk)
         retime_s1_6_reg_reg_IQ <= n_183;
 assign n_159 = retime_s1_6_reg_reg_IQ;
 reg retime_s1_14_reg_reg_IQ;
 always @(posedge clk)
         retime_s1_14_reg_reg_IQ <= n_182;
 assign n_164 = retime_s1_14_reg_reg_IQ;
 reg retime_s1_5_reg_reg_IQ;
 always @(posedge clk)
         retime_s1_5_reg_reg_IQ <= n_185;
 assign n_158 = retime_s1_5_reg_reg_IQ;
 reg retime_s1_3_reg_reg_IQ;
 always @(posedge clk)
         retime_s1_3_reg_reg_IQ <= n_181;
 assign n_156 = retime_s1_3_reg_reg_IQ;
 reg retime_s1_4_reg_reg_IQ;
 always @(posedge clk)
         retime_s1_4_reg_reg_IQ <= n_184;
 assign n_157 = retime_s1_4_reg_reg_IQ;
 reg retime_s1_8_reg_reg_IQ;
 always @(posedge clk)
         retime_s1_8_reg_reg_IQ <= in2_22_0_;
 assign n_27 = retime_s1_8_reg_reg_IQ;
 reg retime_s1_17_reg_reg_IQ;
 always @(posedge clk)
         retime_s1_17_reg_reg_IQ <= {in1[2]};
 assign n_167 = retime_s1_17_reg_reg_IQ;
 reg retime_s1_22_reg_reg_IQ;
 always @(posedge clk)
         retime_s1_22_reg_reg_IQ <= {in2[3]};
 assign n_171 = retime_s1_22_reg_reg_IQ;
 reg retime_s1_21_reg_reg_IQ;
 always @(posedge clk)
         retime_s1_21_reg_reg_IQ <= n_180;
 assign n_25 = retime_s1_21_reg_reg_IQ;
 reg retime_s1_16_reg_reg_IQ;
 always @(posedge clk)
         retime_s1_16_reg_reg_IQ <= {in2[5]};
 assign n_26 = retime_s1_16_reg_reg_IQ;
 reg retime_s1_10_reg_reg_IQ;
 always @(posedge clk)
         retime_s1_10_reg_reg_IQ <= {in1[1]};
 assign n_162 = retime_s1_10_reg_reg_IQ;
 reg retime_s1_20_reg_reg_IQ;
 always @(posedge clk)
         retime_s1_20_reg_reg_IQ <= {in1[5]};
 assign n_169 = retime_s1_20_reg_reg_IQ;
 reg retime_s1_1_reg_reg_IQ;
 always @(posedge clk)
         retime_s1_1_reg_reg_IQ <= {in1[6]};
 assign n_154 = retime_s1_1_reg_reg_IQ;
 reg retime_s1_7_reg_reg_IQ;
 always @(posedge clk)
         retime_s1_7_reg_reg_IQ <= {in1[0]};
 assign n_160 = retime_s1_7_reg_reg_IQ;
 reg retime_s1_11_reg_reg_IQ;
 always @(posedge clk)
         retime_s1_11_reg_reg_IQ <= {in1[3]};
 assign n_163 = retime_s1_11_reg_reg_IQ;
 reg retime_s1_19_reg_reg_IQ;
 always @(posedge clk)
         retime_s1_19_reg_reg_IQ <= {in1[4]};
 assign n_168 = retime_s1_19_reg_reg_IQ;
 reg retime_s1_26_reg_reg_IQ;
 always @(posedge clk)
         retime_s1_26_reg_reg_IQ <= {in2[2]};
 assign n_173 = retime_s1_26_reg_reg_IQ;
 reg retime_s1_15_reg_reg_IQ;
 always @(posedge clk)
         retime_s1_15_reg_reg_IQ <= {in2[4]};
 assign n_165 = retime_s1_15_reg_reg_IQ;
 reg retime_s1_23_reg_reg_IQ;
 always @(posedge clk)
         retime_s1_23_reg_reg_IQ <= {in2[1]};
 assign n_172 = retime_s1_23_reg_reg_IQ;
 reg sub_206_2_retime_s1_9_reg_reg_IQ;
 always @(posedge clk)
         sub_206_2_retime_s1_9_reg_reg_IQ <= sub_206_2_n_79;
 assign sub_206_2_n_85 = sub_206_2_retime_s1_9_reg_reg_IQ;
 reg sub_206_2_retime_s1_25_reg_reg_IQ;
 always @(posedge clk)
         sub_206_2_retime_s1_25_reg_reg_IQ <= in2_20_6_;
 assign sub_206_2_n_81 = sub_206_2_retime_s1_25_reg_reg_IQ;
 reg sub_206_2_retime_s1_13_reg_reg_IQ;
 always @(posedge clk)
         sub_206_2_retime_s1_13_reg_reg_IQ <= sub_206_2_n_77;
 assign sub_206_2_n_83 = sub_206_2_retime_s1_13_reg_reg_IQ;
 reg sub_206_2_retime_s1_18_reg_reg_IQ;
 always @(posedge clk)
         sub_206_2_retime_s1_18_reg_reg_IQ <= sub_206_2_n_78;
 assign sub_206_2_n_82 = sub_206_2_retime_s1_18_reg_reg_IQ;
 reg sub_206_2_retime_s1_12_reg_reg_IQ;
 always @(posedge clk)
         sub_206_2_retime_s1_12_reg_reg_IQ <= {in1[3]};
 assign sub_206_2_n_84 = sub_206_2_retime_s1_12_reg_reg_IQ;
 reg sub_309_2_retime_s1_24_reg_reg_IQ;
 always @(posedge clk)
         sub_309_2_retime_s1_24_reg_reg_IQ <= sub_309_2_n_0;
 assign sub_309_2_n_47 = sub_309_2_retime_s1_24_reg_reg_IQ;
 assign in2_26_6_ = ((in2_25_6_ & ~in2_25_7_) | (in2_23_5_ & in2_25_7_));
 assign in2_26_3_ = ((in2_25_3_ & ~in2_25_7_) | (in2_23_2_ & in2_25_7_));
 assign in2_26_4_ = ((in2_25_4_ & ~in2_25_7_) | (in2_23_3_ & in2_25_7_));
 assign in2_26_5_ = ((in2_25_5_ & ~in2_25_7_) | (in2_23_4_ & in2_25_7_));
 assign in2_26_2_ = ((in2_25_2_ & ~in2_25_7_) | (in2_23_1_ & in2_25_7_));
 assign in2_26_1_ = ((in2_25_1_ & ~in2_25_7_) | (in2_23_0_ & in2_25_7_));
 assign in2_20_6_ = ((in2_19_6_ & ~in2_19_7_) | (in2_17_5_ & in2_19_7_));
 assign in2_29_6_ = ((in2_28_6_ & ~in2_28_7_) | (in2_26_5_ & in2_28_7_));
 assign in2_29_3_ = ((in2_28_3_ & ~in2_28_7_) | (in2_26_2_ & in2_28_7_));
 assign in2_29_4_ = ((in2_28_4_ & ~in2_28_7_) | (in2_26_3_ & in2_28_7_));
 assign in2_29_5_ = ((in2_28_5_ & ~in2_28_7_) | (in2_26_4_ & in2_28_7_));
 assign in2_29_2_ = ((in2_28_2_ & ~in2_28_7_) | (in2_26_1_ & in2_28_7_));
 assign in2_29_1_ = ((in2_28_1_ & ~in2_28_7_) | (in2_26_0_ & in2_28_7_));
 assign in2_17_5_ = ((in2_16_5_ & ~in2_16_7_) | (in2_14_4_ & in2_16_7_));
 assign in2_17_2_ = ((in2_16_2_ & ~in2_16_7_) | (in2_14_1_ & in2_16_7_));
 assign in2_17_1_ = ((in2_16_1_ & ~in2_16_7_) | (in2_14_0_ & in2_16_7_));
 assign in2_17_4_ = ((in2_16_4_ & ~in2_16_7_) | (in2_14_3_ & in2_16_7_));
 assign in2_17_3_ = ((in2_16_3_ & ~in2_16_7_) | (in2_14_2_ & in2_16_7_));
 assign in2_17_0_ = ((in2_16_0_ & ~in2_16_7_) | ({in2[7]} & in2_16_7_));
 assign in2_32_6_ = ((in2_31_6_ & ~in2_31_7_) | (in2_29_5_ & in2_31_7_));
 assign in2_32_3_ = ((in2_31_3_ & ~in2_31_7_) | (in2_29_2_ & in2_31_7_));
 assign in2_32_4_ = ((in2_31_4_ & ~in2_31_7_) | (in2_29_3_ & in2_31_7_));
 assign in2_32_5_ = ((in2_31_5_ & ~in2_31_7_) | (in2_29_4_ & in2_31_7_));
 assign in2_32_2_ = ((in2_31_2_ & ~in2_31_7_) | (in2_29_1_ & in2_31_7_));
 assign in2_32_1_ = ((in2_31_1_ & ~in2_31_7_) | (in2_29_0_ & in2_31_7_));
 assign in2_14_4_ = ((in2_13_4_ & ~in2_13_7_) | (in2_11_3_ & in2_13_7_));
 assign in2_14_1_ = ((in2_13_1_ & ~in2_13_7_) | (in2_11_0_ & in2_13_7_));
 assign in2_14_0_ = ((in2_13_0_ & ~in2_13_7_) | ({in2[8]} & in2_13_7_));
 assign in2_14_3_ = ((in2_13_3_ & ~in2_13_7_) | (in2_11_2_ & in2_13_7_));
 assign in2_14_2_ = ((in2_13_2_ & ~in2_13_7_) | (in2_11_1_ & in2_13_7_));
 assign in2_35_6_ = ((in2_34_6_ & ~in2_34_7_) | (in2_32_5_ & in2_34_7_));
 assign in2_35_3_ = ((in2_34_3_ & ~in2_34_7_) | (in2_32_2_ & in2_34_7_));
 assign in2_35_4_ = ((in2_34_4_ & ~in2_34_7_) | (in2_32_3_ & in2_34_7_));
 assign in2_35_5_ = ((in2_34_5_ & ~in2_34_7_) | (in2_32_4_ & in2_34_7_));
 assign in2_35_2_ = ((in2_34_2_ & ~in2_34_7_) | (in2_32_1_ & in2_34_7_));
 assign in2_35_1_ = ((in2_34_1_ & ~in2_34_7_) | (in2_32_0_ & in2_34_7_));
 assign asc001_0_5_ = ~in2_22_7_;
 assign asc001_0_0_ = ~in2_37_7_;
 assign asc001_0_1_ = ~in2_34_7_;
 assign asc001_0_2_ = ~in2_31_7_;
 assign asc001_0_3_ = ~in2_28_7_;
 assign asc001_0_4_ = ~in2_25_7_;
 assign in2_11_3_ = ((in2_10_3_ & ~in2_10_7_) | (in2_8_2_ & in2_10_7_));
 assign in2_11_0_ = ((in2_10_0_ & ~in2_10_7_) | ({in2[9]} & in2_10_7_));
 assign in2_11_2_ = ((in2_10_2_ & ~in2_10_7_) | (in2_8_1_ & in2_10_7_));
 assign in2_11_1_ = ((in2_10_1_ & ~in2_10_7_) | (in2_8_0_ & in2_10_7_));
 assign in2_8_2_ = ((in2_7_2_ & ~in2_7_7_) | (in2_5_1_ & in2_7_7_));
 assign in2_8_1_ = ((in2_7_1_ & ~in2_7_7_) | (in2_5_0_ & in2_7_7_));
 assign in2_8_0_ = ((in2_7_0_ & ~in2_7_7_) | ({in2[10]} & in2_7_7_));
 assign in2_5_1_ = ((in2_4_1_ & ~in2_4_7_) | (in2_2_0_ & in2_4_7_));
 assign in2_5_0_ = ((in2_4_0_ & ~in2_4_7_) | ({in2[11]} & in2_4_7_));
 assign in2_2_0_ = ((in2_1_0_ & ~in2_1_7_) | ({in2[12]} & in2_1_7_));
 assign n_148 = ~asc001_0_3_;
 assign n_149 = ~asc001_0_5_;
 assign n_150 = ~asc001_0_2_;
 assign n_151 = ~asc001_0_0_;
 assign n_152 = ~asc001_0_4_;
 assign n_153 = ~asc001_0_1_;
 assign in2_23_6_ = ((in2_22_6_ & ~in2_22_7_) | (n_158 & in2_22_7_));
 assign in2_23_5_ = ((in2_22_5_ & ~in2_22_7_) | (n_157 & in2_22_7_));
 assign in2_23_4_ = ((in2_22_4_ & ~in2_22_7_) | (n_164 & in2_22_7_));
 assign in2_23_3_ = ((in2_22_3_ & ~in2_22_7_) | (n_155 & in2_22_7_));
 assign in2_23_2_ = ((in2_22_2_ & ~in2_22_7_) | (n_159 & in2_22_7_));
 assign in2_23_1_ = ((in2_22_1_ & ~in2_22_7_) | (n_156 & in2_22_7_));
 assign in2_29_0_ = ((in2_28_0_ & ~in2_28_7_) | (n_171 & in2_28_7_));
 assign in2_32_0_ = ((in2_31_0_ & ~in2_31_7_) | (n_173 & in2_31_7_));
 assign in2_35_0_ = ((in2_34_0_ & ~in2_34_7_) | (n_172 & in2_34_7_));
 assign in2_23_0_ = ((n_27 & ~in2_22_7_) | (n_26 & in2_22_7_));
 assign in2_26_0_ = ((in2_25_0_ & ~in2_25_7_) | (n_165 & in2_25_7_));
 assign n_54 = ~(n_25 | n_150);
 assign n_52 = ~(n_25 | n_152);
 assign n_53 = ~(n_25 | n_148);
 assign n_51 = ~(n_25 | n_149);
 assign n_55 = ~(n_25 | n_153);
 assign n_56 = ~(n_25 | n_151);
 assign n_186 = ((in2_19_2_ & ~in2_19_7_) | (in2_17_1_ & in2_19_7_));
 assign n_185 = ((in2_19_5_ & ~in2_19_7_) | (in2_17_4_ & in2_19_7_));
 assign n_184 = ((in2_19_4_ & ~in2_19_7_) | (in2_17_3_ & in2_19_7_));
 assign n_183 = ((in2_19_1_ & ~in2_19_7_) | (in2_17_0_ & in2_19_7_));
 assign n_182 = ((in2_19_3_ & ~in2_19_7_) | (in2_17_2_ & in2_19_7_));
 assign n_181 = ((in2_19_0_ & ~in2_19_7_) | ({in2[6]} & in2_19_7_));
 assign n_180 = ~rst;
 assign in2_13_7_ = ~((sub_149_2_n_16 & sub_149_2_n_11) | (sub_149_2_n_33 & sub_149_2_n_25));
 assign in2_13_4_ = ~(sub_149_2_n_33 ^ sub_149_2_n_22);
 assign in2_13_3_ = ~(sub_149_2_n_32 ^ sub_149_2_n_21);
 assign sub_149_2_n_33 = ~(sub_149_2_n_30 & sub_149_2_n_26);
 assign sub_149_2_n_32 = ~(sub_149_2_n_29 & sub_149_2_n_9);
 assign in2_13_2_ = ~(sub_149_2_n_27 ^ sub_149_2_n_19);
 assign sub_149_2_n_30 = ~(sub_149_2_n_27 & sub_149_2_n_20);
 assign sub_149_2_n_29 = ~(sub_149_2_n_27 & sub_149_2_n_13);
 assign in2_13_1_ = ~(sub_149_2_n_24 ^ sub_149_2_n_10);
 assign sub_149_2_n_27 = ((in2_11_0_ & sub_149_2_n_10) | ((in2_11_0_ & sub_149_2_n_7) | (sub_149_2_n_7
    & sub_149_2_n_10)));
 assign sub_149_2_n_26 = ~(sub_149_2_n_23 | sub_149_2_n_8);
 assign sub_149_2_n_25 = ~(sub_149_2_n_17 | sub_149_2_n_14);
 assign sub_149_2_n_24 = ~(in2_11_0_ ^ sub_149_2_n_7);
 assign sub_149_2_n_23 = ~(sub_149_2_n_9 | sub_149_2_n_15);
 assign sub_149_2_n_22 = ({in1[4]} ^ in2_11_3_);
 assign sub_149_2_n_21 = ({in1[3]} ^ in2_11_2_);
 assign sub_149_2_n_20 = ~(sub_149_2_n_12 | sub_149_2_n_15);
 assign sub_149_2_n_19 = ~(sub_149_2_n_9 & sub_149_2_n_13);
 assign in2_13_0_ = ({in1[0]} ^ {in2[8]});
 assign sub_149_2_n_17 = ~sub_149_2_n_16;
 assign sub_149_2_n_16 = ~({in1[5]} | {in1[6]});
 assign sub_149_2_n_15 = ~(in2_11_2_ | sub_149_2_n_1);
 assign sub_149_2_n_14 = ~(in2_11_3_ | sub_149_2_n_2);
 assign sub_149_2_n_13 = ~sub_149_2_n_12;
 assign sub_149_2_n_12 = ~(in2_11_1_ | sub_149_2_n_4);
 assign sub_149_2_n_11 = ~({in1[4]} | sub_149_2_n_6);
 assign sub_149_2_n_10 = ~(sub_149_2_n_3 & {in1[0]});
 assign sub_149_2_n_9 = ~(sub_149_2_n_4 & in2_11_1_);
 assign sub_149_2_n_8 = ~({in1[3]} | sub_149_2_n_5);
 assign sub_149_2_n_7 = ~{in1[1]};
 assign sub_149_2_n_6 = ~in2_11_3_;
 assign sub_149_2_n_5 = ~in2_11_2_;
 assign sub_149_2_n_4 = ~{in1[2]};
 assign sub_149_2_n_3 = ~{in2[8]};
 assign sub_149_2_n_2 = ~{in1[4]};
 assign sub_149_2_n_1 = ~{in1[3]};
 assign in2_28_7_ = ~(sub_248_2_n_41 ^ in2_26_6_);
 assign in2_28_6_ = ~(sub_248_2_n_40 ^ sub_248_2_n_22);
 assign in2_28_5_ = ~(sub_248_2_n_39 ^ sub_248_2_n_19);
 assign sub_248_2_n_41 = ~(sub_248_2_n_35 & sub_248_2_n_32);
 assign sub_248_2_n_40 = ~(sub_248_2_n_36 & sub_248_2_n_28);
 assign sub_248_2_n_39 = ((in2_26_3_ & sub_248_2_n_34) | ((in2_26_3_ & sub_248_2_n_5) | (sub_248_2_n_5
    & sub_248_2_n_34)));
 assign in2_28_4_ = ~(sub_248_2_n_34 ^ sub_248_2_n_18);
 assign in2_28_3_ = ~(sub_248_2_n_33 ^ sub_248_2_n_25);
 assign sub_248_2_n_36 = ~(sub_248_2_n_34 & sub_248_2_n_23);
 assign sub_248_2_n_35 = ~(sub_248_2_n_15 & (sub_248_2_n_12 & (sub_248_2_n_13 & sub_248_2_n_34)));
 assign sub_248_2_n_34 = ~(sub_248_2_n_30 & sub_248_2_n_27);
 assign sub_248_2_n_33 = ((in2_26_1_ & sub_248_2_n_26) | ((in2_26_1_ & sub_248_2_n_3) | (sub_248_2_n_3
    & sub_248_2_n_26)));
 assign sub_248_2_n_32 = ((sub_248_2_n_7 & sub_248_2_n_28) | ((sub_248_2_n_7 & n_154) | (n_154 & sub_248_2_n_28)));
 assign in2_28_2_ = ~(sub_248_2_n_26 ^ sub_248_2_n_21);
 assign sub_248_2_n_30 = ~(sub_248_2_n_26 & sub_248_2_n_24);
 assign in2_28_1_ = ~(sub_248_2_n_20 ^ sub_248_2_n_14);
 assign sub_248_2_n_28 = ((sub_248_2_n_6 & sub_248_2_n_11) | ((sub_248_2_n_6 & n_169) | (n_169 & sub_248_2_n_11)));
 assign sub_248_2_n_27 = ((n_163 | sub_248_2_n_0) & (sub_248_2_n_16 | sub_248_2_n_10));
 assign sub_248_2_n_26 = ((in2_26_0_ & sub_248_2_n_14) | ((in2_26_0_ & sub_248_2_n_4) | (sub_248_2_n_4
    & sub_248_2_n_14)));
 assign sub_248_2_n_25 = (n_163 ^ in2_26_2_);
 assign sub_248_2_n_24 = ((in2_26_2_ | sub_248_2_n_2) & (in2_26_1_ | sub_248_2_n_3));
 assign sub_248_2_n_23 = ((in2_26_4_ | sub_248_2_n_8) & (in2_26_3_ | sub_248_2_n_5));
 assign sub_248_2_n_22 = (n_154 ^ in2_26_5_);
 assign sub_248_2_n_21 = ~(in2_26_1_ ^ sub_248_2_n_3);
 assign sub_248_2_n_20 = ~(in2_26_0_ ^ sub_248_2_n_4);
 assign sub_248_2_n_19 = ~(in2_26_4_ ^ sub_248_2_n_8);
 assign sub_248_2_n_18 = ~(in2_26_3_ ^ sub_248_2_n_5);
 assign in2_28_0_ = (n_160 ^ n_171);
 assign sub_248_2_n_16 = ~(sub_248_2_n_3 & in2_26_1_);
 assign sub_248_2_n_15 = ~(sub_248_2_n_9 & n_168);
 assign sub_248_2_n_14 = ~(sub_248_2_n_1 & n_160);
 assign sub_248_2_n_13 = ~(sub_248_2_n_7 & n_154);
 assign sub_248_2_n_12 = ~(sub_248_2_n_6 & n_169);
 assign sub_248_2_n_11 = ~(sub_248_2_n_5 & in2_26_3_);
 assign sub_248_2_n_10 = ~(in2_26_2_ | sub_248_2_n_2);
 assign sub_248_2_n_9 = ~in2_26_3_;
 assign sub_248_2_n_8 = ~n_169;
 assign sub_248_2_n_7 = ~in2_26_5_;
 assign sub_248_2_n_6 = ~in2_26_4_;
 assign sub_248_2_n_5 = ~n_168;
 assign sub_248_2_n_4 = ~n_162;
 assign sub_248_2_n_3 = ~n_167;
 assign sub_248_2_n_2 = ~n_163;
 assign sub_248_2_n_1 = ~n_171;
 assign sub_248_2_n_0 = ~in2_26_2_;
 assign in2_16_5_ = ~(sub_168_2_n_43 ^ sub_168_2_n_24);
 assign in2_16_7_ = ~(sub_168_2_n_39 | sub_168_2_n_34);
 assign sub_168_2_n_43 = ~(sub_168_2_n_40 & sub_168_2_n_16);
 assign in2_16_4_ = ~(sub_168_2_n_38 ^ sub_168_2_n_22);
 assign in2_16_3_ = ~(sub_168_2_n_36 ^ sub_168_2_n_21);
 assign sub_168_2_n_40 = ~(sub_168_2_n_38 & sub_168_2_n_18);
 assign sub_168_2_n_39 = ~(sub_168_2_n_17 | (sub_168_2_n_15 | ({in1[6]} | sub_168_2_n_37)));
 assign sub_168_2_n_37 = ~sub_168_2_n_38;
 assign sub_168_2_n_38 = ~(sub_168_2_n_33 & sub_168_2_n_29);
 assign sub_168_2_n_36 = ~(sub_168_2_n_32 & sub_168_2_n_10);
 assign in2_16_2_ = ~(sub_168_2_n_28 ^ sub_168_2_n_26);
 assign sub_168_2_n_34 = ~(sub_168_2_n_30 | {in1[6]});
 assign sub_168_2_n_33 = ~(sub_168_2_n_28 & sub_168_2_n_20);
 assign sub_168_2_n_32 = ~(sub_168_2_n_28 & sub_168_2_n_13);
 assign in2_16_1_ = ~(sub_168_2_n_23 ^ sub_168_2_n_14);
 assign sub_168_2_n_30 = ~(sub_168_2_n_27 | sub_168_2_n_9);
 assign sub_168_2_n_29 = ~(sub_168_2_n_25 | sub_168_2_n_11);
 assign sub_168_2_n_28 = ((in2_14_0_ & sub_168_2_n_14) | ((in2_14_0_ & sub_168_2_n_5) | (sub_168_2_n_5
    & sub_168_2_n_14)));
 assign sub_168_2_n_27 = ~(sub_168_2_n_16 | sub_168_2_n_15);
 assign sub_168_2_n_26 = ~(sub_168_2_n_10 & sub_168_2_n_13);
 assign sub_168_2_n_25 = ~(sub_168_2_n_10 | sub_168_2_n_8);
 assign sub_168_2_n_24 = ({in1[5]} ^ in2_14_4_);
 assign sub_168_2_n_23 = ~(in2_14_0_ ^ sub_168_2_n_5);
 assign sub_168_2_n_22 = ~(sub_168_2_n_16 & sub_168_2_n_18);
 assign sub_168_2_n_21 = ({in1[3]} ^ in2_14_2_);
 assign sub_168_2_n_20 = ~(sub_168_2_n_12 | sub_168_2_n_8);
 assign in2_16_0_ = ({in1[0]} ^ {in2[7]});
 assign sub_168_2_n_18 = ~sub_168_2_n_17;
 assign sub_168_2_n_17 = ~(in2_14_3_ | sub_168_2_n_0);
 assign sub_168_2_n_16 = ~(sub_168_2_n_0 & in2_14_3_);
 assign sub_168_2_n_15 = ~(in2_14_4_ | sub_168_2_n_6);
 assign sub_168_2_n_14 = ~(sub_168_2_n_1 & {in1[0]});
 assign sub_168_2_n_13 = ~sub_168_2_n_12;
 assign sub_168_2_n_12 = ~(in2_14_1_ | sub_168_2_n_4);
 assign sub_168_2_n_11 = ~({in1[3]} | sub_168_2_n_3);
 assign sub_168_2_n_10 = ~(sub_168_2_n_4 & in2_14_1_);
 assign sub_168_2_n_9 = ~({in1[5]} | sub_168_2_n_2);
 assign sub_168_2_n_8 = ~(in2_14_2_ | sub_168_2_n_7);
 assign sub_168_2_n_7 = ~{in1[3]};
 assign sub_168_2_n_6 = ~{in1[5]};
 assign sub_168_2_n_5 = ~{in1[1]};
 assign sub_168_2_n_4 = ~{in1[2]};
 assign sub_168_2_n_3 = ~in2_14_2_;
 assign sub_168_2_n_2 = ~in2_14_4_;
 assign sub_168_2_n_1 = ~{in2[7]};
 assign sub_168_2_n_0 = ~{in1[4]};
 assign in2_19_6_ = ~(sub_187_2_n_55 ^ sub_187_2_n_31);
 assign in2_19_5_ = ~(sub_187_2_n_54 ^ sub_187_2_n_30);
 assign in2_19_7_ = ~(sub_187_2_n_49 | sub_187_2_n_46);
 assign sub_187_2_n_55 = ~(sub_187_2_n_51 & sub_187_2_n_38);
 assign sub_187_2_n_54 = ~(sub_187_2_n_50 & sub_187_2_n_22);
 assign in2_19_4_ = ~(sub_187_2_n_47 ^ sub_187_2_n_27);
 assign in2_19_3_ = ~(sub_187_2_n_45 ^ sub_187_2_n_25);
 assign sub_187_2_n_51 = ~(sub_187_2_n_47 & sub_187_2_n_35);
 assign sub_187_2_n_50 = ~(sub_187_2_n_47 & sub_187_2_n_23);
 assign sub_187_2_n_49 = ~sub_187_2_n_48;
 assign sub_187_2_n_48 = ~(sub_187_2_n_23 & (sub_187_2_n_13 & (sub_187_2_n_11 & sub_187_2_n_47)));
 assign sub_187_2_n_47 = ~(sub_187_2_n_41 & sub_187_2_n_36);
 assign sub_187_2_n_46 = ~(sub_187_2_n_43 & sub_187_2_n_18);
 assign sub_187_2_n_45 = ~(sub_187_2_n_42 & sub_187_2_n_15);
 assign in2_19_2_ = ~(sub_187_2_n_37 ^ sub_187_2_n_26);
 assign sub_187_2_n_43 = ~(sub_187_2_n_39 & sub_187_2_n_11);
 assign sub_187_2_n_42 = ~(sub_187_2_n_37 & sub_187_2_n_17);
 assign sub_187_2_n_41 = ~(sub_187_2_n_37 & sub_187_2_n_34);
 assign in2_19_1_ = ~(sub_187_2_n_24 ^ sub_187_2_n_21);
 assign sub_187_2_n_39 = ~sub_187_2_n_38;
 assign sub_187_2_n_38 = ~(sub_187_2_n_33 | sub_187_2_n_20);
 assign sub_187_2_n_37 = ((in2_17_0_ & sub_187_2_n_21) | ((in2_17_0_ & sub_187_2_n_5) | (sub_187_2_n_5
    & sub_187_2_n_21)));
 assign sub_187_2_n_36 = ~(sub_187_2_n_29 | sub_187_2_n_19);
 assign sub_187_2_n_35 = ~sub_187_2_n_32;
 assign sub_187_2_n_34 = ~(sub_187_2_n_16 | sub_187_2_n_14);
 assign sub_187_2_n_33 = ~(sub_187_2_n_22 | sub_187_2_n_12);
 assign sub_187_2_n_32 = ~(sub_187_2_n_23 & sub_187_2_n_13);
 assign sub_187_2_n_31 = ~(sub_187_2_n_18 & sub_187_2_n_11);
 assign sub_187_2_n_30 = ({in1[5]} ^ in2_17_4_);
 assign sub_187_2_n_29 = ~(sub_187_2_n_15 | sub_187_2_n_14);
 assign in2_19_0_ = ({in1[0]} ^ {in2[6]});
 assign sub_187_2_n_27 = ~(sub_187_2_n_22 & sub_187_2_n_23);
 assign sub_187_2_n_26 = ~(sub_187_2_n_15 & sub_187_2_n_17);
 assign sub_187_2_n_25 = ({in1[3]} ^ in2_17_2_);
 assign sub_187_2_n_24 = ~(in2_17_0_ ^ sub_187_2_n_5);
 assign sub_187_2_n_20 = ~({in1[5]} | sub_187_2_n_8);
 assign sub_187_2_n_19 = ~({in1[3]} | sub_187_2_n_6);
 assign sub_187_2_n_23 = ~(sub_187_2_n_0 & {in1[4]});
 assign sub_187_2_n_22 = ~(sub_187_2_n_3 & in2_17_3_);
 assign sub_187_2_n_21 = ~(sub_187_2_n_4 & {in1[0]});
 assign sub_187_2_n_17 = ~sub_187_2_n_16;
 assign sub_187_2_n_13 = ~sub_187_2_n_12;
 assign sub_187_2_n_18 = ~(sub_187_2_n_1 & in2_17_5_);
 assign sub_187_2_n_16 = ~(in2_17_1_ | sub_187_2_n_10);
 assign sub_187_2_n_15 = ~(sub_187_2_n_10 & in2_17_1_);
 assign sub_187_2_n_14 = ~(in2_17_2_ | sub_187_2_n_2);
 assign sub_187_2_n_12 = ~(in2_17_4_ | sub_187_2_n_7);
 assign sub_187_2_n_11 = ~(sub_187_2_n_9 & {in1[6]});
 assign sub_187_2_n_10 = ~{in1[2]};
 assign sub_187_2_n_9 = ~in2_17_5_;
 assign sub_187_2_n_8 = ~in2_17_4_;
 assign sub_187_2_n_7 = ~{in1[5]};
 assign sub_187_2_n_6 = ~in2_17_2_;
 assign sub_187_2_n_5 = ~{in1[1]};
 assign sub_187_2_n_4 = ~{in2[6]};
 assign sub_187_2_n_3 = ~{in1[4]};
 assign sub_187_2_n_2 = ~{in1[3]};
 assign sub_187_2_n_1 = ~{in1[6]};
 assign sub_187_2_n_0 = ~in2_17_3_;
 assign in2_31_7_ = ~(sub_269_2_n_41 ^ in2_29_6_);
 assign in2_31_6_ = ~(sub_269_2_n_40 ^ sub_269_2_n_22);
 assign in2_31_5_ = ~(sub_269_2_n_39 ^ sub_269_2_n_19);
 assign sub_269_2_n_41 = ~(sub_269_2_n_35 & sub_269_2_n_32);
 assign sub_269_2_n_40 = ~(sub_269_2_n_36 & sub_269_2_n_28);
 assign sub_269_2_n_39 = ((in2_29_3_ & sub_269_2_n_34) | ((in2_29_3_ & sub_269_2_n_5) | (sub_269_2_n_5
    & sub_269_2_n_34)));
 assign in2_31_4_ = ~(sub_269_2_n_34 ^ sub_269_2_n_18);
 assign in2_31_3_ = ~(sub_269_2_n_33 ^ sub_269_2_n_25);
 assign sub_269_2_n_36 = ~(sub_269_2_n_34 & sub_269_2_n_23);
 assign sub_269_2_n_35 = ~(sub_269_2_n_15 & (sub_269_2_n_12 & (sub_269_2_n_13 & sub_269_2_n_34)));
 assign sub_269_2_n_34 = ~(sub_269_2_n_30 & sub_269_2_n_27);
 assign sub_269_2_n_33 = ((in2_29_1_ & sub_269_2_n_26) | ((in2_29_1_ & sub_269_2_n_3) | (sub_269_2_n_3
    & sub_269_2_n_26)));
 assign sub_269_2_n_32 = ((sub_269_2_n_7 & sub_269_2_n_28) | ((sub_269_2_n_7 & n_154) | (n_154 & sub_269_2_n_28)));
 assign in2_31_2_ = ~(sub_269_2_n_26 ^ sub_269_2_n_21);
 assign sub_269_2_n_30 = ~(sub_269_2_n_26 & sub_269_2_n_24);
 assign in2_31_1_ = ~(sub_269_2_n_20 ^ sub_269_2_n_14);
 assign sub_269_2_n_28 = ((sub_269_2_n_6 & sub_269_2_n_11) | ((sub_269_2_n_6 & n_169) | (n_169 & sub_269_2_n_11)));
 assign sub_269_2_n_27 = ((n_163 | sub_269_2_n_0) & (sub_269_2_n_16 | sub_269_2_n_10));
 assign sub_269_2_n_26 = ((in2_29_0_ & sub_269_2_n_14) | ((in2_29_0_ & sub_269_2_n_4) | (sub_269_2_n_4
    & sub_269_2_n_14)));
 assign sub_269_2_n_25 = (n_163 ^ in2_29_2_);
 assign sub_269_2_n_24 = ((in2_29_2_ | sub_269_2_n_2) & (in2_29_1_ | sub_269_2_n_3));
 assign sub_269_2_n_23 = ((in2_29_4_ | sub_269_2_n_8) & (in2_29_3_ | sub_269_2_n_5));
 assign sub_269_2_n_22 = (n_154 ^ in2_29_5_);
 assign sub_269_2_n_21 = ~(in2_29_1_ ^ sub_269_2_n_3);
 assign sub_269_2_n_20 = ~(in2_29_0_ ^ sub_269_2_n_4);
 assign sub_269_2_n_19 = ~(in2_29_4_ ^ sub_269_2_n_8);
 assign sub_269_2_n_18 = ~(in2_29_3_ ^ sub_269_2_n_5);
 assign in2_31_0_ = (n_160 ^ n_173);
 assign sub_269_2_n_16 = ~(sub_269_2_n_3 & in2_29_1_);
 assign sub_269_2_n_15 = ~(sub_269_2_n_9 & n_168);
 assign sub_269_2_n_14 = ~(sub_269_2_n_1 & n_160);
 assign sub_269_2_n_13 = ~(sub_269_2_n_7 & n_154);
 assign sub_269_2_n_12 = ~(sub_269_2_n_6 & n_169);
 assign sub_269_2_n_11 = ~(sub_269_2_n_5 & in2_29_3_);
 assign sub_269_2_n_10 = ~(in2_29_2_ | sub_269_2_n_2);
 assign sub_269_2_n_9 = ~in2_29_3_;
 assign sub_269_2_n_8 = ~n_169;
 assign sub_269_2_n_7 = ~in2_29_5_;
 assign sub_269_2_n_6 = ~in2_29_4_;
 assign sub_269_2_n_5 = ~n_168;
 assign sub_269_2_n_4 = ~n_162;
 assign sub_269_2_n_3 = ~n_167;
 assign sub_269_2_n_2 = ~n_163;
 assign sub_269_2_n_1 = ~n_173;
 assign sub_269_2_n_0 = ~in2_29_2_;
 assign in2_34_7_ = ~(sub_290_2_n_41 ^ in2_32_6_);
 assign in2_34_6_ = ~(sub_290_2_n_40 ^ sub_290_2_n_22);
 assign in2_34_5_ = ~(sub_290_2_n_39 ^ sub_290_2_n_19);
 assign sub_290_2_n_41 = ~(sub_290_2_n_35 & sub_290_2_n_32);
 assign sub_290_2_n_40 = ~(sub_290_2_n_36 & sub_290_2_n_28);
 assign sub_290_2_n_39 = ((in2_32_3_ & sub_290_2_n_34) | ((in2_32_3_ & sub_290_2_n_5) | (sub_290_2_n_5
    & sub_290_2_n_34)));
 assign in2_34_4_ = ~(sub_290_2_n_34 ^ sub_290_2_n_18);
 assign in2_34_3_ = ~(sub_290_2_n_33 ^ sub_290_2_n_25);
 assign sub_290_2_n_36 = ~(sub_290_2_n_34 & sub_290_2_n_23);
 assign sub_290_2_n_35 = ~(sub_290_2_n_15 & (sub_290_2_n_12 & (sub_290_2_n_13 & sub_290_2_n_34)));
 assign sub_290_2_n_34 = ~(sub_290_2_n_30 & sub_290_2_n_27);
 assign sub_290_2_n_33 = ((in2_32_1_ & sub_290_2_n_26) | ((in2_32_1_ & sub_290_2_n_3) | (sub_290_2_n_3
    & sub_290_2_n_26)));
 assign sub_290_2_n_32 = ((sub_290_2_n_7 & sub_290_2_n_28) | ((sub_290_2_n_7 & n_154) | (n_154 & sub_290_2_n_28)));
 assign in2_34_2_ = ~(sub_290_2_n_26 ^ sub_290_2_n_21);
 assign sub_290_2_n_30 = ~(sub_290_2_n_26 & sub_290_2_n_24);
 assign in2_34_1_ = ~(sub_290_2_n_20 ^ sub_290_2_n_14);
 assign sub_290_2_n_28 = ((sub_290_2_n_6 & sub_290_2_n_11) | ((sub_290_2_n_6 & n_169) | (n_169 & sub_290_2_n_11)));
 assign sub_290_2_n_27 = ((n_163 | sub_290_2_n_0) & (sub_290_2_n_16 | sub_290_2_n_10));
 assign sub_290_2_n_26 = ((in2_32_0_ & sub_290_2_n_14) | ((in2_32_0_ & sub_290_2_n_4) | (sub_290_2_n_4
    & sub_290_2_n_14)));
 assign sub_290_2_n_25 = (n_163 ^ in2_32_2_);
 assign sub_290_2_n_24 = ((in2_32_2_ | sub_290_2_n_2) & (in2_32_1_ | sub_290_2_n_3));
 assign sub_290_2_n_23 = ((in2_32_4_ | sub_290_2_n_8) & (in2_32_3_ | sub_290_2_n_5));
 assign sub_290_2_n_22 = (n_154 ^ in2_32_5_);
 assign sub_290_2_n_21 = ~(in2_32_1_ ^ sub_290_2_n_3);
 assign sub_290_2_n_20 = ~(in2_32_0_ ^ sub_290_2_n_4);
 assign sub_290_2_n_19 = ~(in2_32_4_ ^ sub_290_2_n_8);
 assign sub_290_2_n_18 = ~(in2_32_3_ ^ sub_290_2_n_5);
 assign in2_34_0_ = (n_160 ^ n_172);
 assign sub_290_2_n_16 = ~(sub_290_2_n_3 & in2_32_1_);
 assign sub_290_2_n_15 = ~(sub_290_2_n_9 & n_168);
 assign sub_290_2_n_14 = ~(sub_290_2_n_1 & n_160);
 assign sub_290_2_n_13 = ~(sub_290_2_n_7 & n_154);
 assign sub_290_2_n_12 = ~(sub_290_2_n_6 & n_169);
 assign sub_290_2_n_11 = ~(sub_290_2_n_5 & in2_32_3_);
 assign sub_290_2_n_10 = ~(in2_32_2_ | sub_290_2_n_2);
 assign sub_290_2_n_9 = ~in2_32_3_;
 assign sub_290_2_n_8 = ~n_169;
 assign sub_290_2_n_7 = ~in2_32_5_;
 assign sub_290_2_n_6 = ~in2_32_4_;
 assign sub_290_2_n_5 = ~n_168;
 assign sub_290_2_n_4 = ~n_162;
 assign sub_290_2_n_3 = ~n_167;
 assign sub_290_2_n_2 = ~n_163;
 assign sub_290_2_n_1 = ~n_172;
 assign sub_290_2_n_0 = ~in2_32_2_;
 assign in2_22_6_ = ~(sub_206_2_n_48 ^ sub_206_2_n_28);
 assign in2_22_5_ = ~(sub_206_2_n_47 ^ sub_206_2_n_25);
 assign sub_206_2_n_49 = ~(sub_206_2_n_42 & sub_206_2_n_39);
 assign sub_206_2_n_48 = ~(sub_206_2_n_44 & sub_206_2_n_33);
 assign sub_206_2_n_47 = ~(sub_206_2_n_43 & sub_206_2_n_13);
 assign in2_22_4_ = ~(sub_206_2_n_41 ^ sub_206_2_n_24);
 assign in2_22_3_ = ~(sub_206_2_n_40 ^ sub_206_2_n_30);
 assign sub_206_2_n_44 = ~(sub_206_2_n_41 & sub_206_2_n_0);
 assign sub_206_2_n_43 = ~(sub_206_2_n_41 & sub_206_2_n_21);
 assign sub_206_2_n_42 = ~(sub_206_2_n_21 & (sub_206_2_n_17 & (sub_206_2_n_19 & sub_206_2_n_41)));
 assign sub_206_2_n_41 = ~(sub_206_2_n_37 & sub_206_2_n_32);
 assign sub_206_2_n_40 = ~(sub_206_2_n_36 & sub_206_2_n_22);
 assign sub_206_2_n_39 = ~(sub_206_2_n_35 | sub_206_2_n_14);
 assign in2_22_2_ = ~(sub_206_2_n_31 ^ sub_206_2_n_27);
 assign sub_206_2_n_37 = ~(sub_206_2_n_31 & sub_206_2_n_29);
 assign sub_206_2_n_36 = ~(sub_206_2_n_31 & sub_206_2_n_16);
 assign sub_206_2_n_35 = ~(sub_206_2_n_33 | sub_206_2_n_18);
 assign sub_206_2_n_33 = ((sub_206_2_n_8 & sub_206_2_n_13) | ((sub_206_2_n_8 & n_169) | (n_169 & sub_206_2_n_13)));
 assign sub_206_2_n_29 = ~(sub_206_2_n_15 | sub_206_2_n_12);
 assign sub_206_2_n_28 = (n_154 ^ n_158);
 assign sub_206_2_n_27 = ~(sub_206_2_n_22 & sub_206_2_n_16);
 assign sub_206_2_n_26 = ~(n_156 ^ sub_206_2_n_6);
 assign sub_206_2_n_25 = (n_169 ^ n_157);
 assign sub_206_2_n_24 = ~(sub_206_2_n_13 & sub_206_2_n_21);
 assign in2_22_0_ = ({in1[0]} ^ {in2[5]});
 assign sub_206_2_n_21 = ~(sub_206_2_n_11 & n_168);
 assign sub_206_2_n_19 = ~sub_206_2_n_18;
 assign sub_206_2_n_18 = ~(n_158 | sub_206_2_n_10);
 assign sub_206_2_n_17 = ~(sub_206_2_n_8 & n_169);
 assign sub_206_2_n_16 = ~sub_206_2_n_15;
 assign sub_206_2_n_14 = ~(n_154 | sub_206_2_n_9);
 assign sub_206_2_n_13 = ~(sub_206_2_n_7 & n_164);
 assign sub_206_2_n_11 = ~n_164;
 assign sub_206_2_n_10 = ~n_154;
 assign sub_206_2_n_9 = ~n_158;
 assign sub_206_2_n_8 = ~n_157;
 assign sub_206_2_n_7 = ~n_168;
 assign sub_206_2_n_6 = ~n_162;
 assign sub_206_2_n_3 = ~{in2[5]};
 assign sub_206_2_n_2 = ~n_155;
 assign sub_206_2_n_0 = ~sub_206_2_n_1;
 assign sub_206_2_n_1 = ~(sub_206_2_n_21 & sub_206_2_n_17);
 assign sub_206_2_n_31 = ((sub_206_2_n_85 & n_156) | ((sub_206_2_n_85 & sub_206_2_n_6) | (sub_206_2_n_6
    & n_156)));
 assign sub_206_2_n_32 = ((sub_206_2_n_84 | sub_206_2_n_2) & (sub_206_2_n_12 | sub_206_2_n_22));
 assign in2_22_1_ = ~(sub_206_2_n_85 ^ sub_206_2_n_26);
 assign in2_22_7_ = ~(sub_206_2_n_81 ^ sub_206_2_n_49);
 assign sub_206_2_n_30 = (sub_206_2_n_84 ^ n_155);
 assign sub_206_2_n_12 = ~(sub_206_2_n_83 | n_155);
 assign sub_206_2_n_15 = ~(sub_206_2_n_82 | n_159);
 assign sub_206_2_n_22 = ~(sub_206_2_n_82 & n_159);
 assign sub_206_2_n_79 = ~({in1[0]} & sub_206_2_n_3);
 assign sub_206_2_n_78 = ~{in1[2]};
 assign sub_206_2_n_77 = ~{in1[3]};
 assign in2_1_7_ = ~sub_73_2_n_6;
 assign sub_73_2_n_6 = ~({in1[4]} | ({in1[5]} | ({in1[6]} | sub_73_2_n_5)));
 assign sub_73_2_n_5 = ~sub_73_2_n_4;
 assign sub_73_2_n_4 = ~(sub_73_2_n_2 | ({in1[1]} | ({in1[2]} | {in1[3]})));
 assign in2_1_0_ = ({in1[0]} ^ {in2[12]});
 assign sub_73_2_n_2 = ~({in2[12]} | sub_73_2_n_1);
 assign sub_73_2_n_1 = ~{in1[0]};
 assign in2_4_7_ = ~(sub_92_2_n_9 & (sub_92_2_n_5 & (sub_92_2_n_6 & sub_92_2_n_3)));
 assign in2_4_1_ = ~(sub_92_2_n_8 ^ sub_92_2_n_4);
 assign sub_92_2_n_9 = ((in2_2_0_ & sub_92_2_n_4) | ((in2_2_0_ & sub_92_2_n_1) | (sub_92_2_n_1 & sub_92_2_n_4)));
 assign sub_92_2_n_8 = ~(in2_2_0_ ^ sub_92_2_n_1);
 assign in2_4_0_ = ({in1[0]} ^ {in2[11]});
 assign sub_92_2_n_6 = ~({in1[4]} | {in1[5]});
 assign sub_92_2_n_5 = ~({in1[2]} | {in1[3]});
 assign sub_92_2_n_4 = ~(sub_92_2_n_2 & {in1[0]});
 assign sub_92_2_n_3 = ~{in1[6]};
 assign sub_92_2_n_2 = ~{in2[11]};
 assign sub_92_2_n_1 = ~{in1[1]};
 assign in2_7_7_ = ~sub_111_2_n_17;
 assign sub_111_2_n_17 = ~({in1[4]} | ({in1[5]} | ({in1[6]} | sub_111_2_n_16)));
 assign sub_111_2_n_16 = ~((sub_111_2_n_7 & sub_111_2_n_4) | (sub_111_2_n_13 & sub_111_2_n_12));
 assign in2_7_2_ = ~(sub_111_2_n_13 ^ sub_111_2_n_10);
 assign in2_7_1_ = ~(sub_111_2_n_11 ^ sub_111_2_n_6);
 assign sub_111_2_n_13 = ((in2_5_0_ & sub_111_2_n_6) | ((in2_5_0_ & sub_111_2_n_3) | (sub_111_2_n_3 &
    sub_111_2_n_6)));
 assign sub_111_2_n_12 = ~(sub_111_2_n_8 | {in1[3]});
 assign sub_111_2_n_11 = ~(in2_5_0_ ^ sub_111_2_n_3);
 assign sub_111_2_n_10 = ({in1[2]} ^ in2_5_1_);
 assign in2_7_0_ = ({in1[0]} ^ {in2[10]});
 assign sub_111_2_n_8 = ~(in2_5_1_ | sub_111_2_n_5);
 assign sub_111_2_n_7 = ~({in1[2]} | sub_111_2_n_2);
 assign sub_111_2_n_6 = ~(sub_111_2_n_1 & {in1[0]});
 assign sub_111_2_n_5 = ~{in1[2]};
 assign sub_111_2_n_4 = ~{in1[3]};
 assign sub_111_2_n_3 = ~{in1[1]};
 assign sub_111_2_n_2 = ~in2_5_1_;
 assign sub_111_2_n_1 = ~{in2[10]};
 assign in2_25_7_ = ~(sub_227_2_n_41 ^ in2_23_6_);
 assign in2_25_6_ = ~(sub_227_2_n_40 ^ sub_227_2_n_22);
 assign in2_25_5_ = ~(sub_227_2_n_39 ^ sub_227_2_n_19);
 assign sub_227_2_n_41 = ~(sub_227_2_n_35 & sub_227_2_n_32);
 assign sub_227_2_n_40 = ~(sub_227_2_n_36 & sub_227_2_n_28);
 assign sub_227_2_n_39 = ((in2_23_3_ & sub_227_2_n_34) | ((in2_23_3_ & sub_227_2_n_5) | (sub_227_2_n_5
    & sub_227_2_n_34)));
 assign in2_25_4_ = ~(sub_227_2_n_34 ^ sub_227_2_n_18);
 assign in2_25_3_ = ~(sub_227_2_n_33 ^ sub_227_2_n_25);
 assign sub_227_2_n_36 = ~(sub_227_2_n_34 & sub_227_2_n_23);
 assign sub_227_2_n_35 = ~(sub_227_2_n_15 & (sub_227_2_n_12 & (sub_227_2_n_13 & sub_227_2_n_34)));
 assign sub_227_2_n_34 = ~(sub_227_2_n_30 & sub_227_2_n_27);
 assign sub_227_2_n_33 = ((in2_23_1_ & sub_227_2_n_26) | ((in2_23_1_ & sub_227_2_n_3) | (sub_227_2_n_3
    & sub_227_2_n_26)));
 assign sub_227_2_n_32 = ((sub_227_2_n_7 & sub_227_2_n_28) | ((sub_227_2_n_7 & n_154) | (n_154 & sub_227_2_n_28)));
 assign in2_25_2_ = ~(sub_227_2_n_26 ^ sub_227_2_n_21);
 assign sub_227_2_n_30 = ~(sub_227_2_n_26 & sub_227_2_n_24);
 assign in2_25_1_ = ~(sub_227_2_n_20 ^ sub_227_2_n_14);
 assign sub_227_2_n_28 = ((sub_227_2_n_6 & sub_227_2_n_11) | ((sub_227_2_n_6 & n_169) | (n_169 & sub_227_2_n_11)));
 assign sub_227_2_n_27 = ((n_163 | sub_227_2_n_0) & (sub_227_2_n_16 | sub_227_2_n_10));
 assign sub_227_2_n_26 = ((in2_23_0_ & sub_227_2_n_14) | ((in2_23_0_ & sub_227_2_n_4) | (sub_227_2_n_4
    & sub_227_2_n_14)));
 assign sub_227_2_n_25 = (n_163 ^ in2_23_2_);
 assign sub_227_2_n_24 = ((in2_23_2_ | sub_227_2_n_2) & (in2_23_1_ | sub_227_2_n_3));
 assign sub_227_2_n_23 = ((in2_23_4_ | sub_227_2_n_8) & (in2_23_3_ | sub_227_2_n_5));
 assign sub_227_2_n_22 = (n_154 ^ in2_23_5_);
 assign sub_227_2_n_21 = ~(in2_23_1_ ^ sub_227_2_n_3);
 assign sub_227_2_n_20 = ~(in2_23_0_ ^ sub_227_2_n_4);
 assign sub_227_2_n_19 = ~(in2_23_4_ ^ sub_227_2_n_8);
 assign sub_227_2_n_18 = ~(sub_227_2_n_11 & sub_227_2_n_15);
 assign in2_25_0_ = (n_160 ^ n_165);
 assign sub_227_2_n_16 = ~(sub_227_2_n_3 & in2_23_1_);
 assign sub_227_2_n_15 = ~(sub_227_2_n_9 & n_168);
 assign sub_227_2_n_14 = ~(sub_227_2_n_1 & n_160);
 assign sub_227_2_n_13 = ~(sub_227_2_n_7 & n_154);
 assign sub_227_2_n_12 = ~(sub_227_2_n_6 & n_169);
 assign sub_227_2_n_11 = ~(sub_227_2_n_5 & in2_23_3_);
 assign sub_227_2_n_10 = ~(in2_23_2_ | sub_227_2_n_2);
 assign sub_227_2_n_9 = ~in2_23_3_;
 assign sub_227_2_n_8 = ~n_169;
 assign sub_227_2_n_7 = ~in2_23_5_;
 assign sub_227_2_n_6 = ~in2_23_4_;
 assign sub_227_2_n_5 = ~n_168;
 assign sub_227_2_n_4 = ~n_162;
 assign sub_227_2_n_3 = ~n_167;
 assign sub_227_2_n_2 = ~n_163;
 assign sub_227_2_n_1 = ~n_165;
 assign sub_227_2_n_0 = ~in2_23_2_;
 assign in2_37_7_ = ~(sub_309_2_n_25 ^ in2_35_6_);
 assign sub_309_2_n_25 = ~(sub_309_2_n_24 & sub_309_2_n_22);
 assign sub_309_2_n_24 = ~(sub_309_2_n_12 & (sub_309_2_n_14 & (sub_309_2_n_13 & sub_309_2_n_23)));
 assign sub_309_2_n_23 = ~(sub_309_2_n_21 & sub_309_2_n_18);
 assign sub_309_2_n_22 = ((sub_309_2_n_4 & sub_309_2_n_19) | ((sub_309_2_n_4 & n_154) | (n_154 & sub_309_2_n_19)));
 assign sub_309_2_n_21 = ~(sub_309_2_n_20 & sub_309_2_n_17);
 assign sub_309_2_n_19 = ((sub_309_2_n_5 & sub_309_2_n_15) | ((sub_309_2_n_5 & n_169) | (n_169 & sub_309_2_n_15)));
 assign sub_309_2_n_18 = ((n_163 | sub_309_2_n_2) & (sub_309_2_n_16 | sub_309_2_n_10));
 assign sub_309_2_n_17 = ((in2_35_2_ | sub_309_2_n_3) & (in2_35_1_ | sub_309_2_n_8));
 assign sub_309_2_n_16 = ~(sub_309_2_n_8 & in2_35_1_);
 assign sub_309_2_n_15 = ~(sub_309_2_n_1 & in2_35_3_);
 assign sub_309_2_n_14 = ~(sub_309_2_n_5 & n_169);
 assign sub_309_2_n_13 = ~(sub_309_2_n_4 & n_154);
 assign sub_309_2_n_12 = ~(sub_309_2_n_6 & n_168);
 assign sub_309_2_n_10 = ~(in2_35_2_ | sub_309_2_n_3);
 assign sub_309_2_n_9 = ~{in2[0]};
 assign sub_309_2_n_8 = ~n_167;
 assign sub_309_2_n_7 = ~n_162;
 assign sub_309_2_n_6 = ~in2_35_3_;
 assign sub_309_2_n_5 = ~in2_35_4_;
 assign sub_309_2_n_4 = ~in2_35_5_;
 assign sub_309_2_n_3 = ~n_163;
 assign sub_309_2_n_2 = ~in2_35_2_;
 assign sub_309_2_n_1 = ~n_168;
 assign sub_309_2_n_20 = ((sub_309_2_n_47 & sub_309_2_n_7) | ((sub_309_2_n_47 & in2_35_0_) | (in2_35_0_
    & sub_309_2_n_7)));
 assign sub_309_2_n_0 = ~({in1[0]} & sub_309_2_n_9);
 assign in2_10_3_ = ~(sub_130_2_n_25 ^ sub_130_2_n_17);
 assign in2_10_7_ = ~sub_130_2_n_27;
 assign sub_130_2_n_27 = ~({in1[4]} | ({in1[5]} | ({in1[6]} | sub_130_2_n_26)));
 assign sub_130_2_n_26 = ~(sub_130_2_n_23 | sub_130_2_n_20);
 assign sub_130_2_n_25 = ~(sub_130_2_n_22 & sub_130_2_n_7);
 assign in2_10_2_ = ~(sub_130_2_n_19 ^ sub_130_2_n_15);
 assign sub_130_2_n_23 = ~(sub_130_2_n_18 | sub_130_2_n_16);
 assign sub_130_2_n_22 = ~(sub_130_2_n_19 & sub_130_2_n_11);
 assign in2_10_1_ = ~(sub_130_2_n_13 ^ sub_130_2_n_9);
 assign sub_130_2_n_20 = ~(sub_130_2_n_14 & sub_130_2_n_10);
 assign sub_130_2_n_18 = ~sub_130_2_n_19;
 assign sub_130_2_n_19 = ((in2_8_0_ & sub_130_2_n_9) | ((in2_8_0_ & sub_130_2_n_4) | (sub_130_2_n_4 &
    sub_130_2_n_9)));
 assign sub_130_2_n_17 = ~(sub_130_2_n_10 & sub_130_2_n_8);
 assign sub_130_2_n_16 = ~(sub_130_2_n_11 & sub_130_2_n_8);
 assign sub_130_2_n_15 = ~(sub_130_2_n_7 & sub_130_2_n_11);
 assign sub_130_2_n_14 = ~(sub_130_2_n_6 & sub_130_2_n_8);
 assign sub_130_2_n_13 = ~(in2_8_0_ ^ sub_130_2_n_4);
 assign in2_10_0_ = ({in1[0]} ^ {in2[9]});
 assign sub_130_2_n_11 = ~(sub_130_2_n_2 & {in1[2]});
 assign sub_130_2_n_10 = ~(sub_130_2_n_3 & in2_8_2_);
 assign sub_130_2_n_9 = ~(sub_130_2_n_1 & {in1[0]});
 assign sub_130_2_n_8 = ~(sub_130_2_n_5 & {in1[3]});
 assign sub_130_2_n_7 = ~sub_130_2_n_6;
 assign sub_130_2_n_6 = ~({in1[2]} | sub_130_2_n_2);
 assign sub_130_2_n_5 = ~in2_8_2_;
 assign sub_130_2_n_4 = ~{in1[1]};
 assign sub_130_2_n_3 = ~{in1[3]};
 assign sub_130_2_n_2 = ~in2_8_1_;
 assign sub_130_2_n_1 = ~{in2[9]};
endmodule
